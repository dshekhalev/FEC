//
// Project       : PLS DVB-S2
// Author        : Shekhalev Denis (des00)
// Workfile      : dvb_pls_dec_constants.svh
// Description   : DVB PLS decoder constants
//

  //------------------------------------------------------------------------------------------------------
  // Gmatrix define
  //------------------------------------------------------------------------------------------------------

  // matrix in reverse form & reverse row order
  localparam bit [0 : 31] cGMATRIX [6] = '{
    32'b11111111111111111111111111111111,
    32'b00000000000000001111111111111111,
    32'b00000000111111110000000011111111,
    32'b00001111000011110000111100001111,
    32'b00110011001100110011001100110011,
    32'b01010101010101010101010101010101
  };

  //------------------------------------------------------------------------------------------------------
  // PLS scrambler
  //------------------------------------------------------------------------------------------------------

  localparam bit [0 : 63] cSCRAMBLE_WORD = 64'b0111000110011101100000111100100101010011010000100010110111111010;

  //------------------------------------------------------------------------------------------------------
  // Hadamard 32 matrix
  //------------------------------------------------------------------------------------------------------

  localparam bit [31 : 0] cHADAMARD32 [32] = '{
    32'b11111111111111111111111111111111,
    32'b10101010101010101010101010101010,
    32'b11001100110011001100110011001100,
    32'b10011001100110011001100110011001,
    32'b11110000111100001111000011110000,
    32'b10100101101001011010010110100101,
    32'b11000011110000111100001111000011,
    32'b10010110100101101001011010010110,
    32'b11111111000000001111111100000000,
    32'b10101010010101011010101001010101,
    32'b11001100001100111100110000110011,
    32'b10011001011001101001100101100110,
    32'b11110000000011111111000000001111,
    32'b10100101010110101010010101011010,
    32'b11000011001111001100001100111100,
    32'b10010110011010011001011001101001,
    32'b11111111111111110000000000000000,
    32'b10101010101010100101010101010101,
    32'b11001100110011000011001100110011,
    32'b10011001100110010110011001100110,
    32'b11110000111100000000111100001111,
    32'b10100101101001010101101001011010,
    32'b11000011110000110011110000111100,
    32'b10010110100101100110100101101001,
    32'b11111111000000000000000011111111,
    32'b10101010010101010101010110101010,
    32'b11001100001100110011001111001100,
    32'b10011001011001100110011010011001,
    32'b11110000000011110000111111110000,
    32'b10100101010110100101101010100101,
    32'b11000011001111000011110011000011,
    32'b10010110011010010110100110010110
  };

