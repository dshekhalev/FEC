//
// Project       : ldpc 3gpp TS 38.212 v15.7.0
// Author        : Shekhalev Denis (des00)
// Workfile      : ldpc_3gpp_constants.svh
// Description   : 3GPP LDPC codec constants, types, functions
//

  typedef logic [2 : 0] idxLs_t;  // 0...7
  typedef logic [2 : 0] idxZc_t;  // 0...7
  typedef logic [5 : 0] code_t;   // graph1/graph2 [4:46]/[4:42]

  //------------------------------------------------------------------------------------------------------
  // code context for variable decoder
  //------------------------------------------------------------------------------------------------------

  typedef struct packed {
    logic   idxGr;       // graph 1/2
    idxLs_t idxLs;       // 0...7
    idxZc_t idxZc;       // 0...7 use only Zc multiply by pDAT_W
    code_t  code;        // graph1/graph2 [4:46]/[4:42]
    logic   do_punct;    // do 3GPP puncture (1)
  } code_ctx_t;

  //------------------------------------------------------------------------------------------------------
  // Zc[idxLs][idxZc]
  //------------------------------------------------------------------------------------------------------

  localparam int cZC_TAB [8][8]= '{
    // pDAT_W        == 1 pDAT_W        == 1/2  pDAT_W        == 1/2/4  pDAT_W        == 1/2/4/8  -- encoder support
    // pLLR_BY_CYCLE == 1 pLLR_BY_CYCLE == 1/2  pLLR_BY_CYCLE == 1/2/4  pLLR_BY_CYCLE == 1/2/4/8  -- decoder support
    //          0           |          1          |           2          |  3 |  4 |  5 |  6 |   7 |
    '{                    2,                    4,                      8,  16,  32,  64, 128, 256},
    '{ 3,                      6,                    12,                    24,  48,  96, 192, 384}, // | extended |
    '{ 5,                     10,                    20,                    40,  80, 160, 320,              320},
    '{ 7,                     14,                    28,                    56, 112, 224,                   448, 448},
    '{ 9,                     18,                    36,                    72, 144, 288,                   288, 288},
    '{11,                     22,                    44,                    88, 176, 352,                   352, 352},
    '{13,                     26,                    52,                   104, 208,                        416, 416, 416},
    '{15,                     30,                    60,                   120, 240,                        480, 480, 480}
    };

  //------------------------------------------------------------------------------------------------------
  // Main code bit tab [idxGr][idxLs][idxZc][do_punct] == sended data with main LDPC matrix
  //------------------------------------------------------------------------------------------------------

  localparam int cMAIN_CODE_BIT_TAB [2][8][8][2] = '{
    // gr 1
    '{
      '{  '{52, 48},  '{104, 96},  '{208, 192},    '{416, 384},   '{832, 768},   '{1664, 1536},   '{3328, 3072},   '{6656, 6144}},
      '{  '{78, 72}, '{156, 144},  '{312, 288},    '{624, 576}, '{1248, 1152},   '{2496, 2304},   '{4992, 4608},   '{9984, 9216}},
      '{'{130, 120}, '{260, 240},  '{520, 480},   '{1040, 960}, '{2080, 1920},   '{4160, 3840},   '{8320, 7680},   '{8320, 7680}},
      '{'{182, 168}, '{364, 336},  '{728, 672},  '{1456, 1344}, '{2912, 2688},   '{5824, 5376}, '{11648, 10752}, '{11648, 10752}},
      '{'{234, 216}, '{468, 432},  '{936, 864},  '{1872, 1728}, '{3744, 3456},   '{7488, 6912},   '{7488, 6912},   '{7488, 6912}},
      '{'{286, 264}, '{572, 528}, '{1144, 1056}, '{2288, 2112}, '{4576, 4224},   '{9152, 8448},   '{9152, 8448},   '{9152, 8448}},
      '{'{338, 312}, '{676, 624}, '{1352, 1248}, '{2704, 2496}, '{5408, 4992},  '{10816, 9984},  '{10816, 9984},  '{10816, 9984}},
      '{'{390, 360}, '{780, 720}, '{1560, 1440}, '{3120, 2880}, '{6240, 5760}, '{12480, 11520}, '{12480, 11520}, '{12480, 11520}}
    },
    // gr 2
    '{
      '{  '{28, 24},   '{56, 48},  '{112, 96},   '{224, 192},   '{448, 384},   '{896, 768}, '{1792, 1536}, '{3584, 3072}},
      '{  '{42, 36},   '{84, 72}, '{168, 144},   '{336, 288},   '{672, 576}, '{1344, 1152}, '{2688, 2304}, '{5376, 4608}},
      '{  '{70, 60}, '{140, 120}, '{280, 240},   '{560, 480},  '{1120, 960}, '{2240, 1920}, '{4480, 3840}, '{4480, 3840}},
      '{  '{98, 84}, '{196, 168}, '{392, 336},   '{784, 672}, '{1568, 1344}, '{3136, 2688}, '{6272, 5376}, '{6272, 5376}},
      '{'{126, 108}, '{252, 216}, '{504, 432},  '{1008, 864}, '{2016, 1728}, '{4032, 3456}, '{4032, 3456}, '{4032, 3456}},
      '{'{154, 132}, '{308, 264}, '{616, 528}, '{1232, 1056}, '{2464, 2112}, '{4928, 4224}, '{4928, 4224}, '{4928, 4224}},
      '{'{182, 156}, '{364, 312}, '{728, 624}, '{1456, 1248}, '{2912, 2496}, '{5824, 4992}, '{5824, 4992}, '{5824, 4992}},
      '{'{210, 180}, '{420, 360}, '{840, 720}, '{1680, 1440}, '{3360, 2880}, '{6720, 5760}, '{6720, 5760}, '{6720, 5760}}
    }
  };

  //------------------------------------------------------------------------------------------------------
  //
  //------------------------------------------------------------------------------------------------------

  localparam int cZC_MAX        = 480; // 384;
  localparam int cLOG2_ZC_MAX   = 9;

  typedef logic [cLOG2_ZC_MAX-1 : 0] hb_zc_t;

  //------------------------------------------------------------------------------------------------------
  // usefull functions
  //------------------------------------------------------------------------------------------------------

  function automatic int get_data_bit_length (input logic idxGr, idxLs_t idxLs, idxZc_t idxZc);
    if (idxGr) begin
      get_data_bit_length = 10*cZC_TAB[idxLs][idxZc];
    end
    else begin
      get_data_bit_length = 22*cZC_TAB[idxLs][idxZc];
    end
  endfunction

  function automatic int get_code_bit_length (input logic idxGr, idxLs_t idxLs, idxZc_t idxZc, code_t code, logic punct);
    if (code < 4) code = 4;
    //
    if (idxGr) begin
      if (punct) begin
        get_code_bit_length = ( 8 + code)*cZC_TAB[idxLs][idxZc];
      end
      else begin
        get_code_bit_length = (10 + code)*cZC_TAB[idxLs][idxZc];
      end
    end
    else begin
      if (punct) begin
        get_code_bit_length = (20 + code)*cZC_TAB[idxLs][idxZc];
      end
      else begin
        get_code_bit_length = (22 + code)*cZC_TAB[idxLs][idxZc];
      end
    end
  endfunction

  function automatic int get_main_code_bit_length (input logic idxGr, idxLs_t idxLs, idxZc_t idxZc, logic punct);
    get_main_code_bit_length = get_code_bit_length(idxGr, idxLs, idxZc, 4, punct);
  endfunction

  // number of columns for systematic channel LLRs
  localparam int cGR_SYST_BIT_COL   [2] = '{22, 10};

  // number of columns for systematic and major parity channel LLRs
  localparam int cGR_MAJOR_BIT_COL  [2] = '{26, 14};

  // number of maximim rows for whole matix
  localparam int cGR_MAX_ROW        [2] = '{46, 42};

  // number of maximum columns for whole matrix
  localparam int cGR_MAX_COL        [2] = '{68, 52};

  //------------------------------------------------------------------------------------------------------
  // inv(-E*T^-1*B+D) for major check matrix decoder
  //  cINV_PSI[idxGr][idxLs][idxZc]
  //------------------------------------------------------------------------------------------------------

  localparam int cINV_PSI [2][8][8] = '{
    // graph 1
    '{
      '{0, 0, 0, 0,   0, 0, 0, 0},
      '{0, 0, 0, 0,   0, 0, 0, 0},  // | extended |
      '{0, 0, 0, 0,   0, 0, 0,              0},
      '{0, 0, 0, 0,   0, 0,                 0,   0},
      '{0, 0, 0, 0,   0, 0,                 0,   0},
      '{0, 0, 0, 0,   0, 0,                 0,   0},
      '{1, 1, 1, 1, 105,                  105, 105, 105},
      '{0, 0, 0, 0,   0,                    0,   0,   0}
     },
    // graph 2
    '{
      '{1, 1, 1, 1, 1, 1, 1, 1},
      '{1, 1, 1, 1, 1, 1, 1, 1},    // | extended |
      '{1, 1, 1, 1, 1, 1, 1,              1},
      '{0, 0, 0, 0, 0, 0,                 0, 0},
      '{1, 1, 1, 1, 1, 1,                 1, 1},
      '{1, 1, 1, 1, 1, 1,                 1, 1},
      '{1, 1, 1, 1, 1,                    1, 1, 1},
      '{0, 0, 0, 0, 0,                    0, 0, 0}
     }
  };

  //------------------------------------------------------------------------------------------------------
  // check matrix based types
  //------------------------------------------------------------------------------------------------------

  typedef int baseHc_t [46][68];

  typedef logic            [5 : 0] hb_row_t;
  typedef logic            [6 : 0] hb_col_t;
  typedef logic [cLOG2_ZC_MAX : 0] hb_value_t; // {sign, hb_zc_t}

