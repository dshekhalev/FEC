localparam int          cSHORT_HS_TAB_11BY45_PACKED_SIZE = 136;
localparam bit [18 : 0] cSHORT_HS_TAB_11BY45_PACKED[cSHORT_HS_TAB_11BY45_PACKED_SIZE] = '{
{  1'b1, 1'b0,  8'd44,    9'd1},{  1'b0, 1'b0,  8'd11,    9'd0},{  1'b0, 1'b0,   8'd6,   9'd13},{  1'b0, 1'b1,   8'd0,   9'd88},
{  1'b0, 1'b0,  8'd12,    9'd0},{  1'b0, 1'b0,  8'd11,    9'd0},{  1'b0, 1'b0,   8'd8,  9'd311},{  1'b0, 1'b1,   8'd4,  9'd251},
{  1'b0, 1'b0,  8'd13,    9'd0},{  1'b0, 1'b0,  8'd12,    9'd0},{  1'b0, 1'b0,   8'd6,  9'd221},{  1'b0, 1'b1,   8'd4,  9'd247},
{  1'b0, 1'b0,  8'd14,    9'd0},{  1'b0, 1'b0,  8'd13,    9'd0},{  1'b0, 1'b0,  8'd10,   9'd55},{  1'b0, 1'b1,   8'd9,  9'd203},
{  1'b0, 1'b0,  8'd15,    9'd0},{  1'b0, 1'b0,  8'd14,    9'd0},{  1'b0, 1'b0,   8'd4,   9'd94},{  1'b0, 1'b1,   8'd2,   9'd60},
{  1'b0, 1'b0,  8'd16,    9'd0},{  1'b0, 1'b0,  8'd15,    9'd0},{  1'b0, 1'b0,   8'd3,  9'd151},{  1'b0, 1'b1,   8'd0,  9'd217},
{  1'b0, 1'b0,  8'd17,    9'd0},{  1'b0, 1'b0,  8'd16,    9'd0},{  1'b0, 1'b0,   8'd1,   9'd77},{  1'b0, 1'b1,   8'd0,  9'd270},
{  1'b0, 1'b0,  8'd18,    9'd0},{  1'b0, 1'b0,  8'd17,    9'd0},{  1'b0, 1'b0,   8'd3,  9'd249},{  1'b0, 1'b1,   8'd2,  9'd140},
{  1'b0, 1'b0,  8'd19,    9'd0},{  1'b0, 1'b0,  8'd18,    9'd0},{  1'b0, 1'b0,   8'd9,  9'd253},{  1'b0, 1'b1,   8'd8,   9'd42},
{  1'b0, 1'b0,  8'd20,    9'd0},{  1'b0, 1'b0,  8'd19,    9'd0},{  1'b0, 1'b0,   8'd1,  9'd128},{  1'b0, 1'b1,   8'd0,  9'd239},
{  1'b0, 1'b0,  8'd21,    9'd0},{  1'b0, 1'b0,  8'd20,    9'd0},{  1'b0, 1'b0,   8'd2,  9'd166},{  1'b0, 1'b1,   8'd0,  9'd266},
{  1'b0, 1'b0,  8'd22,    9'd0},{  1'b0, 1'b0,  8'd21,    9'd0},{  1'b0, 1'b0,   8'd8,   9'd86},{  1'b0, 1'b1,   8'd7,  9'd337},
{  1'b0, 1'b0,  8'd23,    9'd0},{  1'b0, 1'b0,  8'd22,    9'd0},{  1'b0, 1'b0,   8'd5,  9'd308},{  1'b0, 1'b1,   8'd3,  9'd152},
{  1'b0, 1'b0,  8'd24,    9'd0},{  1'b0, 1'b0,  8'd23,    9'd0},{  1'b0, 1'b0,   8'd2,  9'd104},{  1'b0, 1'b1,   8'd1,  9'd238},
{  1'b0, 1'b0,  8'd25,    9'd0},{  1'b0, 1'b0,  8'd24,    9'd0},{  1'b0, 1'b0,   8'd6,  9'd109},{  1'b0, 1'b1,   8'd0,   9'd29},
{  1'b0, 1'b0,  8'd26,    9'd0},{  1'b0, 1'b0,  8'd25,    9'd0},{  1'b0, 1'b0,   8'd4,   9'd89},{  1'b0, 1'b1,   8'd2,  9'd245},
{  1'b0, 1'b0,  8'd27,    9'd0},{  1'b0, 1'b0,  8'd26,    9'd0},{  1'b0, 1'b0,   8'd7,  9'd323},{  1'b0, 1'b1,   8'd2,   9'd84},
{  1'b0, 1'b0,  8'd28,    9'd0},{  1'b0, 1'b0,  8'd27,    9'd0},{  1'b0, 1'b0,   8'd4,  9'd351},{  1'b0, 1'b1,   8'd0,  9'd357},
{  1'b0, 1'b0,  8'd29,    9'd0},{  1'b0, 1'b0,  8'd28,    9'd0},{  1'b0, 1'b0,   8'd4,   9'd30},{  1'b0, 1'b1,   8'd3,   9'd26},
{  1'b0, 1'b0,  8'd30,    9'd0},{  1'b0, 1'b0,  8'd29,    9'd0},{  1'b0, 1'b0,   8'd3,  9'd148},{  1'b0, 1'b1,   8'd1,  9'd322},
{  1'b0, 1'b0,  8'd31,    9'd0},{  1'b0, 1'b0,  8'd30,    9'd0},{  1'b0, 1'b0,   8'd2,  9'd222},{  1'b0, 1'b1,   8'd1,  9'd324},
{  1'b0, 1'b0,  8'd32,    9'd0},{  1'b0, 1'b0,  8'd31,    9'd0},{  1'b0, 1'b0,   8'd7,   9'd22},{  1'b0, 1'b1,   8'd5,  9'd155},
{  1'b0, 1'b0,  8'd33,    9'd0},{  1'b0, 1'b0,  8'd32,    9'd0},{  1'b0, 1'b0,   8'd3,  9'd281},{  1'b0, 1'b1,   8'd1,  9'd155},
{  1'b0, 1'b0,  8'd34,    9'd0},{  1'b0, 1'b0,  8'd33,    9'd0},{  1'b0, 1'b0,   8'd3,   9'd55},{  1'b0, 1'b1,   8'd1,  9'd271},
{  1'b0, 1'b0,  8'd35,    9'd0},{  1'b0, 1'b0,  8'd34,    9'd0},{  1'b0, 1'b0,  8'd10,  9'd165},{  1'b0, 1'b1,   8'd4,  9'd242},
{  1'b0, 1'b0,  8'd36,    9'd0},{  1'b0, 1'b0,  8'd35,    9'd0},{  1'b0, 1'b0,  8'd10,  9'd187},{  1'b0, 1'b1,   8'd4,   9'd26},
{  1'b0, 1'b0,  8'd37,    9'd0},{  1'b0, 1'b0,  8'd36,    9'd0},{  1'b0, 1'b0,   8'd5,  9'd319},{  1'b0, 1'b1,   8'd3,  9'd237},
{  1'b0, 1'b0,  8'd38,    9'd0},{  1'b0, 1'b0,  8'd37,    9'd0},{  1'b0, 1'b0,   8'd4,  9'd111},{  1'b0, 1'b1,   8'd3,   9'd98},
{  1'b0, 1'b0,  8'd39,    9'd0},{  1'b0, 1'b0,  8'd38,    9'd0},{  1'b0, 1'b0,   8'd2,  9'd352},{  1'b0, 1'b1,   8'd1,  9'd351},
{  1'b0, 1'b0,  8'd40,    9'd0},{  1'b0, 1'b0,  8'd39,    9'd0},{  1'b0, 1'b0,   8'd4,  9'd134},{  1'b0, 1'b1,   8'd2,  9'd257},
{  1'b0, 1'b0,  8'd41,    9'd0},{  1'b0, 1'b0,  8'd40,    9'd0},{  1'b0, 1'b0,   8'd3,  9'd204},{  1'b0, 1'b1,   8'd0,  9'd330},
{  1'b0, 1'b0,  8'd42,    9'd0},{  1'b0, 1'b0,  8'd41,    9'd0},{  1'b0, 1'b0,   8'd9,  9'd331},{  1'b0, 1'b1,   8'd0,  9'd138},
{  1'b0, 1'b0,  8'd43,    9'd0},{  1'b0, 1'b0,  8'd42,    9'd0},{  1'b0, 1'b0,   8'd2,  9'd205},{  1'b0, 1'b1,   8'd1,  9'd359},
{  1'b0, 1'b0,  8'd44,    9'd0},{  1'b0, 1'b0,  8'd43,    9'd0},{  1'b0, 1'b0,   8'd1,  9'd209},{  1'b0, 1'b1,   8'd0,  9'd189}
};
localparam bit [18 : 0] cSHORT_HS_V_TAB_11BY45_PACKED[cSHORT_HS_TAB_11BY45_PACKED_SIZE] = '{
{ 8'd44, 1'b0,   10'd0},{ 8'd44, 1'b1, 10'd132},
{ 8'd43, 1'b0, 10'd128},{ 8'd43, 1'b1, 10'd133},
{ 8'd42, 1'b0, 10'd124},{ 8'd42, 1'b1, 10'd129},
{ 8'd41, 1'b0, 10'd120},{ 8'd41, 1'b1, 10'd125},
{ 8'd40, 1'b0, 10'd116},{ 8'd40, 1'b1, 10'd121},
{ 8'd39, 1'b0, 10'd112},{ 8'd39, 1'b1, 10'd117},
{ 8'd38, 1'b0, 10'd108},{ 8'd38, 1'b1, 10'd113},
{ 8'd37, 1'b0, 10'd104},{ 8'd37, 1'b1, 10'd109},
{ 8'd36, 1'b0, 10'd100},{ 8'd36, 1'b1, 10'd105},
{ 8'd35, 1'b0,  10'd96},{ 8'd35, 1'b1, 10'd101},
{ 8'd34, 1'b0,  10'd92},{ 8'd34, 1'b1,  10'd97},
{ 8'd33, 1'b0,  10'd88},{ 8'd33, 1'b1,  10'd93},
{ 8'd32, 1'b0,  10'd84},{ 8'd32, 1'b1,  10'd89},
{ 8'd31, 1'b0,  10'd80},{ 8'd31, 1'b1,  10'd85},
{ 8'd30, 1'b0,  10'd76},{ 8'd30, 1'b1,  10'd81},
{ 8'd29, 1'b0,  10'd72},{ 8'd29, 1'b1,  10'd77},
{ 8'd28, 1'b0,  10'd68},{ 8'd28, 1'b1,  10'd73},
{ 8'd27, 1'b0,  10'd64},{ 8'd27, 1'b1,  10'd69},
{ 8'd26, 1'b0,  10'd60},{ 8'd26, 1'b1,  10'd65},
{ 8'd25, 1'b0,  10'd56},{ 8'd25, 1'b1,  10'd61},
{ 8'd24, 1'b0,  10'd52},{ 8'd24, 1'b1,  10'd57},
{ 8'd23, 1'b0,  10'd48},{ 8'd23, 1'b1,  10'd53},
{ 8'd22, 1'b0,  10'd44},{ 8'd22, 1'b1,  10'd49},
{ 8'd21, 1'b0,  10'd40},{ 8'd21, 1'b1,  10'd45},
{ 8'd20, 1'b0,  10'd36},{ 8'd20, 1'b1,  10'd41},
{ 8'd19, 1'b0,  10'd32},{ 8'd19, 1'b1,  10'd37},
{ 8'd18, 1'b0,  10'd28},{ 8'd18, 1'b1,  10'd33},
{ 8'd17, 1'b0,  10'd24},{ 8'd17, 1'b1,  10'd29},
{ 8'd16, 1'b0,  10'd20},{ 8'd16, 1'b1,  10'd25},
{ 8'd15, 1'b0,  10'd16},{ 8'd15, 1'b1,  10'd21},
{ 8'd14, 1'b0,  10'd12},{ 8'd14, 1'b1,  10'd17},
{ 8'd13, 1'b0,   10'd8},{ 8'd13, 1'b1,  10'd13},
{ 8'd12, 1'b0,   10'd4},{ 8'd12, 1'b1,   10'd9},
{ 8'd11, 1'b0,   10'd1},{ 8'd11, 1'b1,   10'd5},
{ 8'd10, 1'b0,  10'd14},{ 8'd10, 1'b0,  10'd98},{ 8'd10, 1'b1, 10'd102},
{  8'd9, 1'b0,  10'd15},{  8'd9, 1'b0,  10'd34},{  8'd9, 1'b1, 10'd126},
{  8'd8, 1'b0,   10'd6},{  8'd8, 1'b0,  10'd35},{  8'd8, 1'b1,  10'd46},
{  8'd7, 1'b0,  10'd47},{  8'd7, 1'b0,  10'd66},{  8'd7, 1'b1,  10'd86},
{  8'd6, 1'b0,   10'd2},{  8'd6, 1'b0,  10'd10},{  8'd6, 1'b1,  10'd58},
{  8'd5, 1'b0,  10'd50},{  8'd5, 1'b0,  10'd87},{  8'd5, 1'b1, 10'd106},
{  8'd4, 1'b0,   10'd7},{  8'd4, 1'b0,  10'd11},{  8'd4, 1'b0,  10'd18},{  8'd4, 1'b0,  10'd62},{  8'd4, 1'b0,  10'd70},{  8'd4, 1'b0,  10'd74},{  8'd4, 1'b0,  10'd99},{  8'd4, 1'b0, 10'd103},{  8'd4, 1'b0, 10'd110},{  8'd4, 1'b1, 10'd118},
{  8'd3, 1'b0,  10'd22},{  8'd3, 1'b0,  10'd30},{  8'd3, 1'b0,  10'd51},{  8'd3, 1'b0,  10'd75},{  8'd3, 1'b0,  10'd78},{  8'd3, 1'b0,  10'd90},{  8'd3, 1'b0,  10'd94},{  8'd3, 1'b0, 10'd107},{  8'd3, 1'b0, 10'd111},{  8'd3, 1'b1, 10'd122},
{  8'd2, 1'b0,  10'd19},{  8'd2, 1'b0,  10'd31},{  8'd2, 1'b0,  10'd42},{  8'd2, 1'b0,  10'd54},{  8'd2, 1'b0,  10'd63},{  8'd2, 1'b0,  10'd67},{  8'd2, 1'b0,  10'd82},{  8'd2, 1'b0, 10'd114},{  8'd2, 1'b0, 10'd119},{  8'd2, 1'b1, 10'd130},
{  8'd1, 1'b0,  10'd26},{  8'd1, 1'b0,  10'd38},{  8'd1, 1'b0,  10'd55},{  8'd1, 1'b0,  10'd79},{  8'd1, 1'b0,  10'd83},{  8'd1, 1'b0,  10'd91},{  8'd1, 1'b0,  10'd95},{  8'd1, 1'b0, 10'd115},{  8'd1, 1'b0, 10'd131},{  8'd1, 1'b1, 10'd134},
{  8'd0, 1'b0,   10'd3},{  8'd0, 1'b0,  10'd23},{  8'd0, 1'b0,  10'd27},{  8'd0, 1'b0,  10'd39},{  8'd0, 1'b0,  10'd43},{  8'd0, 1'b0,  10'd59},{  8'd0, 1'b0,  10'd71},{  8'd0, 1'b0, 10'd123},{  8'd0, 1'b0, 10'd127},{  8'd0, 1'b1, 10'd135}
};
localparam int          cSHORT_HS_TAB_4BY15_PACKED_SIZE = 162;
localparam bit [18 : 0] cSHORT_HS_TAB_4BY15_PACKED[cSHORT_HS_TAB_4BY15_PACKED_SIZE] = '{
{  1'b0, 1'b0,  8'd26,    9'd0},{  1'b0, 1'b0,  8'd25,    9'd0},{  1'b0, 1'b0,  8'd10,  9'd354},{  1'b0, 1'b1,   8'd2,   9'd69},
{  1'b0, 1'b0,  8'd32,    9'd0},{  1'b0, 1'b0,  8'd31,    9'd0},{  1'b0, 1'b0,   8'd4,  9'd225},{  1'b0, 1'b1,   8'd2,  9'd270},
{  1'b0, 1'b0,  8'd34,    9'd0},{  1'b0, 1'b0,  8'd33,    9'd0},{  1'b0, 1'b0,   8'd7,  9'd149},{  1'b0, 1'b1,   8'd1,  9'd333},
{  1'b1, 1'b0,  8'd44,    9'd1},{  1'b0, 1'b0,  8'd12,    9'd0},{  1'b0, 1'b0,   8'd6,  9'd356},{  1'b0, 1'b0,   8'd2,  9'd167},{  1'b0, 1'b1,   8'd0,  9'd141},
{  1'b0, 1'b0,  8'd13,    9'd0},{  1'b0, 1'b0,  8'd12,    9'd0},{  1'b0, 1'b0,   8'd8,   9'd69},{  1'b0, 1'b0,   8'd2,  9'd137},{  1'b0, 1'b1,   8'd0,  9'd255},
{  1'b0, 1'b0,  8'd14,    9'd0},{  1'b0, 1'b0,  8'd13,    9'd0},{  1'b0, 1'b0,   8'd5,  9'd261},{  1'b0, 1'b0,   8'd2,  9'd100},{  1'b0, 1'b1,   8'd1,  9'd287},
{  1'b0, 1'b0,  8'd15,    9'd0},{  1'b0, 1'b0,  8'd14,    9'd0},{  1'b0, 1'b0,   8'd6,  9'd243},{  1'b0, 1'b0,   8'd1,  9'd157},{  1'b0, 1'b1,   8'd0,  9'd305},
{  1'b0, 1'b0,  8'd16,    9'd0},{  1'b0, 1'b0,  8'd15,    9'd0},{  1'b0, 1'b0,   8'd8,  9'd113},{  1'b0, 1'b0,   8'd1,  9'd316},{  1'b0, 1'b1,   8'd0,   9'd77},
{  1'b0, 1'b0,  8'd17,    9'd0},{  1'b0, 1'b0,  8'd16,    9'd0},{  1'b0, 1'b0,   8'd3,  9'd302},{  1'b0, 1'b0,   8'd1,  9'd338},{  1'b0, 1'b1,   8'd0,  9'd233},
{  1'b0, 1'b0,  8'd18,    9'd0},{  1'b0, 1'b0,  8'd17,    9'd0},{  1'b0, 1'b0,   8'd9,  9'd136},{  1'b0, 1'b0,   8'd2,  9'd206},{  1'b0, 1'b1,   8'd0,   9'd59},
{  1'b0, 1'b0,  8'd19,    9'd0},{  1'b0, 1'b0,  8'd18,    9'd0},{  1'b0, 1'b0,   8'd5,  9'd206},{  1'b0, 1'b0,   8'd1,  9'd238},{  1'b0, 1'b1,   8'd0,  9'd278},
{  1'b0, 1'b0,  8'd20,    9'd0},{  1'b0, 1'b0,  8'd19,    9'd0},{  1'b0, 1'b0,  8'd10,  9'd334},{  1'b0, 1'b0,   8'd1,  9'd276},{  1'b0, 1'b1,   8'd0,  9'd290},
{  1'b0, 1'b0,  8'd21,    9'd0},{  1'b0, 1'b0,  8'd20,    9'd0},{  1'b0, 1'b0,   8'd3,   9'd59},{  1'b0, 1'b0,   8'd2,  9'd299},{  1'b0, 1'b1,   8'd1,  9'd228},
{  1'b0, 1'b0,  8'd22,    9'd0},{  1'b0, 1'b0,  8'd21,    9'd0},{  1'b0, 1'b0,   8'd8,  9'd303},{  1'b0, 1'b0,   8'd2,  9'd277},{  1'b0, 1'b1,   8'd1,   9'd72},
{  1'b0, 1'b0,  8'd23,    9'd0},{  1'b0, 1'b0,  8'd22,    9'd0},{  1'b0, 1'b0,   8'd3,  9'd273},{  1'b0, 1'b0,   8'd1,  9'd349},{  1'b0, 1'b1,   8'd0,  9'd208},
{  1'b0, 1'b0,  8'd24,    9'd0},{  1'b0, 1'b0,  8'd23,    9'd0},{  1'b0, 1'b0,   8'd7,  9'd353},{  1'b0, 1'b0,   8'd2,  9'd224},{  1'b0, 1'b1,   8'd1,   9'd74},
{  1'b0, 1'b0,  8'd25,    9'd0},{  1'b0, 1'b0,  8'd24,    9'd0},{  1'b0, 1'b0,   8'd4,    9'd0},{  1'b0, 1'b0,   8'd1,   9'd62},{  1'b0, 1'b1,   8'd0,  9'd265},
{  1'b0, 1'b0,  8'd27,    9'd0},{  1'b0, 1'b0,  8'd26,    9'd0},{  1'b0, 1'b0,   8'd3,  9'd229},{  1'b0, 1'b0,   8'd1,  9'd351},{  1'b0, 1'b1,   8'd0,  9'd230},
{  1'b0, 1'b0,  8'd28,    9'd0},{  1'b0, 1'b0,  8'd27,    9'd0},{  1'b0, 1'b0,   8'd7,  9'd316},{  1'b0, 1'b0,   8'd2,   9'd39},{  1'b0, 1'b1,   8'd0,   9'd79},
{  1'b0, 1'b0,  8'd29,    9'd0},{  1'b0, 1'b0,  8'd28,    9'd0},{  1'b0, 1'b0,   8'd7,  9'd268},{  1'b0, 1'b0,   8'd1,   9'd64},{  1'b0, 1'b1,   8'd0,  9'd354},
{  1'b0, 1'b0,  8'd30,    9'd0},{  1'b0, 1'b0,  8'd29,    9'd0},{  1'b0, 1'b0,   8'd6,  9'd303},{  1'b0, 1'b0,   8'd2,  9'd110},{  1'b0, 1'b1,   8'd0,  9'd289},
{  1'b0, 1'b0,  8'd31,    9'd0},{  1'b0, 1'b0,  8'd30,    9'd0},{  1'b0, 1'b0,  8'd11,  9'd317},{  1'b0, 1'b0,   8'd2,   9'd52},{  1'b0, 1'b1,   8'd1,   9'd15},
{  1'b0, 1'b0,  8'd33,    9'd0},{  1'b0, 1'b0,  8'd32,    9'd0},{  1'b0, 1'b0,   8'd9,  9'd241},{  1'b0, 1'b0,   8'd2,   9'd14},{  1'b0, 1'b1,   8'd0,   9'd70},
{  1'b0, 1'b0,  8'd35,    9'd0},{  1'b0, 1'b0,  8'd34,    9'd0},{  1'b0, 1'b0,   8'd9,  9'd322},{  1'b0, 1'b0,   8'd2,  9'd245},{  1'b0, 1'b1,   8'd0,  9'd195},
{  1'b0, 1'b0,  8'd36,    9'd0},{  1'b0, 1'b0,  8'd35,    9'd0},{  1'b0, 1'b0,   8'd4,  9'd253},{  1'b0, 1'b0,   8'd1,  9'd200},{  1'b0, 1'b1,   8'd0,  9'd172},
{  1'b0, 1'b0,  8'd37,    9'd0},{  1'b0, 1'b0,  8'd36,    9'd0},{  1'b0, 1'b0,   8'd5,  9'd338},{  1'b0, 1'b0,   8'd2,  9'd296},{  1'b0, 1'b1,   8'd1,   9'd23},
{  1'b0, 1'b0,  8'd38,    9'd0},{  1'b0, 1'b0,  8'd37,    9'd0},{  1'b0, 1'b0,   8'd5,  9'd207},{  1'b0, 1'b0,   8'd2,  9'd200},{  1'b0, 1'b1,   8'd1,  9'd344},
{  1'b0, 1'b0,  8'd39,    9'd0},{  1'b0, 1'b0,  8'd38,    9'd0},{  1'b0, 1'b0,   8'd4,   9'd47},{  1'b0, 1'b0,   8'd1,  9'd206},{  1'b0, 1'b1,   8'd0,  9'd238},
{  1'b0, 1'b0,  8'd40,    9'd0},{  1'b0, 1'b0,  8'd39,    9'd0},{  1'b0, 1'b0,   8'd8,  9'd189},{  1'b0, 1'b0,   8'd2,  9'd326},{  1'b0, 1'b1,   8'd0,  9'd347},
{  1'b0, 1'b0,  8'd41,    9'd0},{  1'b0, 1'b0,  8'd40,    9'd0},{  1'b0, 1'b0,  8'd11,   9'd94},{  1'b0, 1'b0,   8'd2,  9'd241},{  1'b0, 1'b1,   8'd0,  9'd151},
{  1'b0, 1'b0,  8'd42,    9'd0},{  1'b0, 1'b0,  8'd41,    9'd0},{  1'b0, 1'b0,   8'd6,  9'd241},{  1'b0, 1'b0,   8'd2,  9'd234},{  1'b0, 1'b1,   8'd1,  9'd102},
{  1'b0, 1'b0,  8'd43,    9'd0},{  1'b0, 1'b0,  8'd42,    9'd0},{  1'b0, 1'b0,  8'd11,  9'd301},{  1'b0, 1'b0,   8'd2,  9'd127},{  1'b0, 1'b1,   8'd1,  9'd290},
{  1'b0, 1'b0,  8'd44,    9'd0},{  1'b0, 1'b0,  8'd43,    9'd0},{  1'b0, 1'b0,  8'd10,  9'd269},{  1'b0, 1'b0,   8'd2,  9'd359},{  1'b0, 1'b1,   8'd0,  9'd300}
};
localparam bit [18 : 0] cSHORT_HS_V_TAB_4BY15_PACKED[cSHORT_HS_TAB_4BY15_PACKED_SIZE] = '{
{ 8'd44, 1'b0,  10'd12},{ 8'd44, 1'b1, 10'd157},
{ 8'd43, 1'b0, 10'd152},{ 8'd43, 1'b1, 10'd158},
{ 8'd42, 1'b0, 10'd147},{ 8'd42, 1'b1, 10'd153},
{ 8'd41, 1'b0, 10'd142},{ 8'd41, 1'b1, 10'd148},
{ 8'd40, 1'b0, 10'd137},{ 8'd40, 1'b1, 10'd143},
{ 8'd39, 1'b0, 10'd132},{ 8'd39, 1'b1, 10'd138},
{ 8'd38, 1'b0, 10'd127},{ 8'd38, 1'b1, 10'd133},
{ 8'd37, 1'b0, 10'd122},{ 8'd37, 1'b1, 10'd128},
{ 8'd36, 1'b0, 10'd117},{ 8'd36, 1'b1, 10'd123},
{ 8'd35, 1'b0, 10'd112},{ 8'd35, 1'b1, 10'd118},
{ 8'd34, 1'b0,   10'd8},{ 8'd34, 1'b1, 10'd113},
{ 8'd33, 1'b0, 10'd107},{ 8'd33, 1'b1,   10'd9},
{ 8'd32, 1'b0,   10'd4},{ 8'd32, 1'b1, 10'd108},
{ 8'd31, 1'b0, 10'd102},{ 8'd31, 1'b1,   10'd5},
{ 8'd30, 1'b0,  10'd97},{ 8'd30, 1'b1, 10'd103},
{ 8'd29, 1'b0,  10'd92},{ 8'd29, 1'b1,  10'd98},
{ 8'd28, 1'b0,  10'd87},{ 8'd28, 1'b1,  10'd93},
{ 8'd27, 1'b0,  10'd82},{ 8'd27, 1'b1,  10'd88},
{ 8'd26, 1'b0,   10'd0},{ 8'd26, 1'b1,  10'd83},
{ 8'd25, 1'b0,  10'd77},{ 8'd25, 1'b1,   10'd1},
{ 8'd24, 1'b0,  10'd72},{ 8'd24, 1'b1,  10'd78},
{ 8'd23, 1'b0,  10'd67},{ 8'd23, 1'b1,  10'd73},
{ 8'd22, 1'b0,  10'd62},{ 8'd22, 1'b1,  10'd68},
{ 8'd21, 1'b0,  10'd57},{ 8'd21, 1'b1,  10'd63},
{ 8'd20, 1'b0,  10'd52},{ 8'd20, 1'b1,  10'd58},
{ 8'd19, 1'b0,  10'd47},{ 8'd19, 1'b1,  10'd53},
{ 8'd18, 1'b0,  10'd42},{ 8'd18, 1'b1,  10'd48},
{ 8'd17, 1'b0,  10'd37},{ 8'd17, 1'b1,  10'd43},
{ 8'd16, 1'b0,  10'd32},{ 8'd16, 1'b1,  10'd38},
{ 8'd15, 1'b0,  10'd27},{ 8'd15, 1'b1,  10'd33},
{ 8'd14, 1'b0,  10'd22},{ 8'd14, 1'b1,  10'd28},
{ 8'd13, 1'b0,  10'd17},{ 8'd13, 1'b1,  10'd23},
{ 8'd12, 1'b0,  10'd13},{ 8'd12, 1'b1,  10'd18},
{ 8'd11, 1'b0, 10'd104},{ 8'd11, 1'b0, 10'd144},{ 8'd11, 1'b1, 10'd154},
{ 8'd10, 1'b0,  10'd54},{ 8'd10, 1'b0,   10'd2},{ 8'd10, 1'b1, 10'd159},
{  8'd9, 1'b0,  10'd44},{  8'd9, 1'b0, 10'd109},{  8'd9, 1'b1, 10'd114},
{  8'd8, 1'b0,  10'd19},{  8'd8, 1'b0,  10'd34},{  8'd8, 1'b0,  10'd64},{  8'd8, 1'b1, 10'd139},
{  8'd7, 1'b0,  10'd74},{  8'd7, 1'b0,  10'd89},{  8'd7, 1'b0,  10'd94},{  8'd7, 1'b1,  10'd10},
{  8'd6, 1'b0,  10'd14},{  8'd6, 1'b0,  10'd29},{  8'd6, 1'b0,  10'd99},{  8'd6, 1'b1, 10'd149},
{  8'd5, 1'b0,  10'd24},{  8'd5, 1'b0,  10'd49},{  8'd5, 1'b0, 10'd124},{  8'd5, 1'b1, 10'd129},
{  8'd4, 1'b0,  10'd79},{  8'd4, 1'b0,   10'd6},{  8'd4, 1'b0, 10'd119},{  8'd4, 1'b1, 10'd134},
{  8'd3, 1'b0,  10'd39},{  8'd3, 1'b0,  10'd59},{  8'd3, 1'b0,  10'd69},{  8'd3, 1'b1,  10'd84},
{  8'd2, 1'b0,  10'd15},{  8'd2, 1'b0,  10'd20},{  8'd2, 1'b0,  10'd25},{  8'd2, 1'b0,  10'd45},{  8'd2, 1'b0,  10'd60},{  8'd2, 1'b0,  10'd65},{  8'd2, 1'b0,  10'd75},{  8'd2, 1'b0,   10'd3},{  8'd2, 1'b0,  10'd90},{  8'd2, 1'b0, 10'd100},{  8'd2, 1'b0, 10'd105},{  8'd2, 1'b0,   10'd7},{  8'd2, 1'b0, 10'd110},{  8'd2, 1'b0, 10'd115},{  8'd2, 1'b0, 10'd125},{  8'd2, 1'b0, 10'd130},{  8'd2, 1'b0, 10'd140},{  8'd2, 1'b0, 10'd145},{  8'd2, 1'b0, 10'd150},{  8'd2, 1'b0, 10'd155},{  8'd2, 1'b1, 10'd160},
{  8'd1, 1'b0,  10'd26},{  8'd1, 1'b0,  10'd30},{  8'd1, 1'b0,  10'd35},{  8'd1, 1'b0,  10'd40},{  8'd1, 1'b0,  10'd50},{  8'd1, 1'b0,  10'd55},{  8'd1, 1'b0,  10'd61},{  8'd1, 1'b0,  10'd66},{  8'd1, 1'b0,  10'd70},{  8'd1, 1'b0,  10'd76},{  8'd1, 1'b0,  10'd80},{  8'd1, 1'b0,  10'd85},{  8'd1, 1'b0,  10'd95},{  8'd1, 1'b0, 10'd106},{  8'd1, 1'b0,  10'd11},{  8'd1, 1'b0, 10'd120},{  8'd1, 1'b0, 10'd126},{  8'd1, 1'b0, 10'd131},{  8'd1, 1'b0, 10'd135},{  8'd1, 1'b0, 10'd151},{  8'd1, 1'b1, 10'd156},
{  8'd0, 1'b0,  10'd16},{  8'd0, 1'b0,  10'd21},{  8'd0, 1'b0,  10'd31},{  8'd0, 1'b0,  10'd36},{  8'd0, 1'b0,  10'd41},{  8'd0, 1'b0,  10'd46},{  8'd0, 1'b0,  10'd51},{  8'd0, 1'b0,  10'd56},{  8'd0, 1'b0,  10'd71},{  8'd0, 1'b0,  10'd81},{  8'd0, 1'b0,  10'd86},{  8'd0, 1'b0,  10'd91},{  8'd0, 1'b0,  10'd96},{  8'd0, 1'b0, 10'd101},{  8'd0, 1'b0, 10'd111},{  8'd0, 1'b0, 10'd116},{  8'd0, 1'b0, 10'd121},{  8'd0, 1'b0, 10'd136},{  8'd0, 1'b0, 10'd141},{  8'd0, 1'b0, 10'd146},{  8'd0, 1'b1, 10'd161}
};
localparam int          cSHORT_HS_TAB_14BY45_PACKED_SIZE = 155;
localparam bit [18 : 0] cSHORT_HS_TAB_14BY45_PACKED[cSHORT_HS_TAB_14BY45_PACKED_SIZE] = '{
{  1'b1, 1'b0,  8'd44,    9'd1},{  1'b0, 1'b0,  8'd14,    9'd0},{  1'b0, 1'b0,  8'd11,  9'd310},{  1'b0, 1'b0,   8'd9,  9'd156},{  1'b0, 1'b1,   8'd6,  9'd173},
{  1'b0, 1'b0,  8'd15,    9'd0},{  1'b0, 1'b0,  8'd14,    9'd0},{  1'b0, 1'b0,   8'd4,   9'd19},{  1'b0, 1'b0,   8'd3,  9'd183},{  1'b0, 1'b1,   8'd2,  9'd320},
{  1'b0, 1'b0,  8'd16,    9'd0},{  1'b0, 1'b0,  8'd15,    9'd0},{  1'b0, 1'b0,   8'd3,  9'd263},{  1'b0, 1'b0,   8'd1,  9'd294},{  1'b0, 1'b1,   8'd0,  9'd297},
{  1'b0, 1'b0,  8'd17,    9'd0},{  1'b0, 1'b0,  8'd16,    9'd0},{  1'b0, 1'b0,   8'd3,   9'd45},{  1'b0, 1'b0,   8'd1,  9'd150},{  1'b0, 1'b1,   8'd0,  9'd137},
{  1'b0, 1'b0,  8'd18,    9'd0},{  1'b0, 1'b0,  8'd17,    9'd0},{  1'b0, 1'b0,   8'd4,   9'd95},{  1'b0, 1'b0,   8'd3,  9'd170},{  1'b0, 1'b1,   8'd2,   9'd97},
{  1'b0, 1'b0,  8'd19,    9'd0},{  1'b0, 1'b0,  8'd18,    9'd0},{  1'b0, 1'b0,  8'd13,  9'd105},{  1'b0, 1'b0,   8'd5,   9'd30},{  1'b0, 1'b1,   8'd3,  9'd132},
{  1'b0, 1'b0,  8'd20,    9'd0},{  1'b0, 1'b0,  8'd19,    9'd0},{  1'b0, 1'b0,   8'd3,   9'd85},{  1'b0, 1'b0,   8'd2,   9'd48},{  1'b0, 1'b1,   8'd0,  9'd257},
{  1'b0, 1'b0,  8'd21,    9'd0},{  1'b0, 1'b0,  8'd20,    9'd0},{  1'b0, 1'b0,  8'd10,  9'd125},{  1'b0, 1'b0,   8'd5,   9'd91},{  1'b0, 1'b1,   8'd4,  9'd211},
{  1'b0, 1'b0,  8'd22,    9'd0},{  1'b0, 1'b0,  8'd21,    9'd0},{  1'b0, 1'b0,  8'd12,  9'd359},{  1'b0, 1'b0,   8'd2,   9'd43},{  1'b0, 1'b1,   8'd0,  9'd147},
{  1'b0, 1'b0,  8'd23,    9'd0},{  1'b0, 1'b0,  8'd22,    9'd0},{  1'b0, 1'b0,   8'd9,  9'd218},{  1'b0, 1'b0,   8'd4,   9'd34},{  1'b0, 1'b1,   8'd0,  9'd306},
{  1'b0, 1'b0,  8'd24,    9'd0},{  1'b0, 1'b0,  8'd23,    9'd0},{  1'b0, 1'b0,   8'd6,  9'd230},{  1'b0, 1'b0,   8'd4,    9'd0},{  1'b0, 1'b1,   8'd0,  9'd217},
{  1'b0, 1'b0,  8'd25,    9'd0},{  1'b0, 1'b0,  8'd24,    9'd0},{  1'b0, 1'b0,   8'd5,  9'd205},{  1'b0, 1'b0,   8'd3,  9'd253},{  1'b0, 1'b1,   8'd0,  9'd252},
{  1'b0, 1'b0,  8'd26,    9'd0},{  1'b0, 1'b0,  8'd25,    9'd0},{  1'b0, 1'b0,   8'd8,  9'd172},{  1'b0, 1'b0,   8'd7,  9'd156},{  1'b0, 1'b1,   8'd1,  9'd264},
{  1'b0, 1'b0,  8'd27,    9'd0},{  1'b0, 1'b0,  8'd26,    9'd0},{  1'b0, 1'b0,   8'd4,   9'd20},{  1'b0, 1'b0,   8'd2,  9'd273},{  1'b0, 1'b1,   8'd1,  9'd132},
{  1'b0, 1'b0,  8'd28,    9'd0},{  1'b0, 1'b0,  8'd27,    9'd0},{  1'b0, 1'b0,  8'd12,  9'd203},{  1'b0, 1'b0,  8'd10,  9'd355},{  1'b0, 1'b1,   8'd4,  9'd185},
{  1'b0, 1'b0,  8'd29,    9'd0},{  1'b0, 1'b0,  8'd28,    9'd0},{  1'b0, 1'b0,  8'd11,  9'd132},{  1'b0, 1'b0,   8'd6,  9'd240},{  1'b0, 1'b1,   8'd5,  9'd101},
{  1'b0, 1'b0,  8'd30,    9'd0},{  1'b0, 1'b0,  8'd29,    9'd0},{  1'b0, 1'b0,   8'd5,  9'd245},{  1'b0, 1'b0,   8'd4,   9'd86},{  1'b0, 1'b1,   8'd3,  9'd276},
{  1'b0, 1'b0,  8'd31,    9'd0},{  1'b0, 1'b0,  8'd30,    9'd0},{  1'b0, 1'b0,   8'd7,   9'd15},{  1'b0, 1'b0,   8'd3,  9'd235},{  1'b0, 1'b1,   8'd1,  9'd125},
{  1'b0, 1'b0,  8'd32,    9'd0},{  1'b0, 1'b0,  8'd31,    9'd0},{  1'b0, 1'b0,   8'd4,  9'd184},{  1'b0, 1'b0,   8'd2,  9'd251},{  1'b0, 1'b1,   8'd1,  9'd214},
{  1'b0, 1'b0,  8'd33,    9'd0},{  1'b0, 1'b0,  8'd32,    9'd0},{  1'b0, 1'b0,  8'd12,  9'd139},{  1'b0, 1'b0,   8'd8,   9'd52},{  1'b0, 1'b1,   8'd1,  9'd354},
{  1'b0, 1'b0,  8'd34,    9'd0},{  1'b0, 1'b0,  8'd33,    9'd0},{  1'b0, 1'b0,   8'd4,  9'd195},{  1'b0, 1'b0,   8'd2,  9'd175},{  1'b0, 1'b1,   8'd1,  9'd247},
{  1'b0, 1'b0,  8'd35,    9'd0},{  1'b0, 1'b0,  8'd34,    9'd0},{  1'b0, 1'b0,   8'd4,    9'd6},{  1'b0, 1'b0,   8'd3,  9'd120},{  1'b0, 1'b1,   8'd0,  9'd116},
{  1'b0, 1'b0,  8'd36,    9'd0},{  1'b0, 1'b0,  8'd35,    9'd0},{  1'b0, 1'b0,   8'd5,    9'd2},{  1'b0, 1'b0,   8'd2,  9'd164},{  1'b0, 1'b1,   8'd0,  9'd302},
{  1'b0, 1'b0,  8'd37,    9'd0},{  1'b0, 1'b0,  8'd36,    9'd0},{  1'b0, 1'b0,  8'd13,  9'd254},{  1'b0, 1'b0,   8'd5,  9'd153},{  1'b0, 1'b1,   8'd2,  9'd159},
{  1'b0, 1'b0,  8'd38,    9'd0},{  1'b0, 1'b0,  8'd37,    9'd0},{  1'b0, 1'b0,   8'd2,  9'd204},{  1'b0, 1'b0,   8'd1,   9'd29},{  1'b0, 1'b1,   8'd0,  9'd135},
{  1'b0, 1'b0,  8'd39,    9'd0},{  1'b0, 1'b0,  8'd38,    9'd0},{  1'b0, 1'b0,   8'd9,  9'd184},{  1'b0, 1'b0,   8'd2,   9'd26},{  1'b0, 1'b1,   8'd0,   9'd51},
{  1'b0, 1'b0,  8'd40,    9'd0},{  1'b0, 1'b0,  8'd39,    9'd0},{  1'b0, 1'b0,   8'd8,  9'd272},{  1'b0, 1'b0,   8'd5,    9'd4},{  1'b0, 1'b1,   8'd4,   9'd67},
{  1'b0, 1'b0,  8'd41,    9'd0},{  1'b0, 1'b0,  8'd40,    9'd0},{  1'b0, 1'b0,  8'd13,  9'd122},{  1'b0, 1'b0,   8'd5,   9'd12},{  1'b0, 1'b1,   8'd2,  9'd210},
{  1'b0, 1'b0,  8'd42,    9'd0},{  1'b0, 1'b0,  8'd41,    9'd0},{  1'b0, 1'b0,   8'd7,  9'd299},{  1'b0, 1'b0,   8'd1,  9'd114},{  1'b0, 1'b1,   8'd0,   9'd12},
{  1'b0, 1'b0,  8'd43,    9'd0},{  1'b0, 1'b0,  8'd42,    9'd0},{  1'b0, 1'b0,  8'd11,  9'd175},{  1'b0, 1'b0,   8'd3,  9'd182},{  1'b0, 1'b1,   8'd1,  9'd181},
{  1'b0, 1'b0,  8'd44,    9'd0},{  1'b0, 1'b0,  8'd43,    9'd0},{  1'b0, 1'b0,  8'd10,  9'd143},{  1'b0, 1'b0,   8'd3,  9'd358},{  1'b0, 1'b1,   8'd1,   9'd31}
};
localparam bit [18 : 0] cSHORT_HS_V_TAB_14BY45_PACKED[cSHORT_HS_TAB_14BY45_PACKED_SIZE] = '{
{ 8'd44, 1'b0,   10'd0},{ 8'd44, 1'b1, 10'd150},
{ 8'd43, 1'b0, 10'd145},{ 8'd43, 1'b1, 10'd151},
{ 8'd42, 1'b0, 10'd140},{ 8'd42, 1'b1, 10'd146},
{ 8'd41, 1'b0, 10'd135},{ 8'd41, 1'b1, 10'd141},
{ 8'd40, 1'b0, 10'd130},{ 8'd40, 1'b1, 10'd136},
{ 8'd39, 1'b0, 10'd125},{ 8'd39, 1'b1, 10'd131},
{ 8'd38, 1'b0, 10'd120},{ 8'd38, 1'b1, 10'd126},
{ 8'd37, 1'b0, 10'd115},{ 8'd37, 1'b1, 10'd121},
{ 8'd36, 1'b0, 10'd110},{ 8'd36, 1'b1, 10'd116},
{ 8'd35, 1'b0, 10'd105},{ 8'd35, 1'b1, 10'd111},
{ 8'd34, 1'b0, 10'd100},{ 8'd34, 1'b1, 10'd106},
{ 8'd33, 1'b0,  10'd95},{ 8'd33, 1'b1, 10'd101},
{ 8'd32, 1'b0,  10'd90},{ 8'd32, 1'b1,  10'd96},
{ 8'd31, 1'b0,  10'd85},{ 8'd31, 1'b1,  10'd91},
{ 8'd30, 1'b0,  10'd80},{ 8'd30, 1'b1,  10'd86},
{ 8'd29, 1'b0,  10'd75},{ 8'd29, 1'b1,  10'd81},
{ 8'd28, 1'b0,  10'd70},{ 8'd28, 1'b1,  10'd76},
{ 8'd27, 1'b0,  10'd65},{ 8'd27, 1'b1,  10'd71},
{ 8'd26, 1'b0,  10'd60},{ 8'd26, 1'b1,  10'd66},
{ 8'd25, 1'b0,  10'd55},{ 8'd25, 1'b1,  10'd61},
{ 8'd24, 1'b0,  10'd50},{ 8'd24, 1'b1,  10'd56},
{ 8'd23, 1'b0,  10'd45},{ 8'd23, 1'b1,  10'd51},
{ 8'd22, 1'b0,  10'd40},{ 8'd22, 1'b1,  10'd46},
{ 8'd21, 1'b0,  10'd35},{ 8'd21, 1'b1,  10'd41},
{ 8'd20, 1'b0,  10'd30},{ 8'd20, 1'b1,  10'd36},
{ 8'd19, 1'b0,  10'd25},{ 8'd19, 1'b1,  10'd31},
{ 8'd18, 1'b0,  10'd20},{ 8'd18, 1'b1,  10'd26},
{ 8'd17, 1'b0,  10'd15},{ 8'd17, 1'b1,  10'd21},
{ 8'd16, 1'b0,  10'd10},{ 8'd16, 1'b1,  10'd16},
{ 8'd15, 1'b0,   10'd5},{ 8'd15, 1'b1,  10'd11},
{ 8'd14, 1'b0,   10'd1},{ 8'd14, 1'b1,   10'd6},
{ 8'd13, 1'b0,  10'd27},{ 8'd13, 1'b0, 10'd117},{ 8'd13, 1'b1, 10'd137},
{ 8'd12, 1'b0,  10'd42},{ 8'd12, 1'b0,  10'd72},{ 8'd12, 1'b1,  10'd97},
{ 8'd11, 1'b0,   10'd2},{ 8'd11, 1'b0,  10'd77},{ 8'd11, 1'b1, 10'd147},
{ 8'd10, 1'b0,  10'd37},{ 8'd10, 1'b0,  10'd73},{ 8'd10, 1'b1, 10'd152},
{  8'd9, 1'b0,   10'd3},{  8'd9, 1'b0,  10'd47},{  8'd9, 1'b1, 10'd127},
{  8'd8, 1'b0,  10'd62},{  8'd8, 1'b0,  10'd98},{  8'd8, 1'b1, 10'd132},
{  8'd7, 1'b0,  10'd63},{  8'd7, 1'b0,  10'd87},{  8'd7, 1'b1, 10'd142},
{  8'd6, 1'b0,   10'd4},{  8'd6, 1'b0,  10'd52},{  8'd6, 1'b1,  10'd78},
{  8'd5, 1'b0,  10'd28},{  8'd5, 1'b0,  10'd38},{  8'd5, 1'b0,  10'd57},{  8'd5, 1'b0,  10'd79},{  8'd5, 1'b0,  10'd82},{  8'd5, 1'b0, 10'd112},{  8'd5, 1'b0, 10'd118},{  8'd5, 1'b0, 10'd133},{  8'd5, 1'b1, 10'd138},
{  8'd4, 1'b0,   10'd7},{  8'd4, 1'b0,  10'd22},{  8'd4, 1'b0,  10'd39},{  8'd4, 1'b0,  10'd48},{  8'd4, 1'b0,  10'd53},{  8'd4, 1'b0,  10'd67},{  8'd4, 1'b0,  10'd74},{  8'd4, 1'b0,  10'd83},{  8'd4, 1'b0,  10'd92},{  8'd4, 1'b0, 10'd102},{  8'd4, 1'b0, 10'd107},{  8'd4, 1'b1, 10'd134},
{  8'd3, 1'b0,   10'd8},{  8'd3, 1'b0,  10'd12},{  8'd3, 1'b0,  10'd17},{  8'd3, 1'b0,  10'd23},{  8'd3, 1'b0,  10'd29},{  8'd3, 1'b0,  10'd32},{  8'd3, 1'b0,  10'd58},{  8'd3, 1'b0,  10'd84},{  8'd3, 1'b0,  10'd88},{  8'd3, 1'b0, 10'd108},{  8'd3, 1'b0, 10'd148},{  8'd3, 1'b1, 10'd153},
{  8'd2, 1'b0,   10'd9},{  8'd2, 1'b0,  10'd24},{  8'd2, 1'b0,  10'd33},{  8'd2, 1'b0,  10'd43},{  8'd2, 1'b0,  10'd68},{  8'd2, 1'b0,  10'd93},{  8'd2, 1'b0, 10'd103},{  8'd2, 1'b0, 10'd113},{  8'd2, 1'b0, 10'd119},{  8'd2, 1'b0, 10'd122},{  8'd2, 1'b0, 10'd128},{  8'd2, 1'b1, 10'd139},
{  8'd1, 1'b0,  10'd13},{  8'd1, 1'b0,  10'd18},{  8'd1, 1'b0,  10'd64},{  8'd1, 1'b0,  10'd69},{  8'd1, 1'b0,  10'd89},{  8'd1, 1'b0,  10'd94},{  8'd1, 1'b0,  10'd99},{  8'd1, 1'b0, 10'd104},{  8'd1, 1'b0, 10'd123},{  8'd1, 1'b0, 10'd143},{  8'd1, 1'b0, 10'd149},{  8'd1, 1'b1, 10'd154},
{  8'd0, 1'b0,  10'd14},{  8'd0, 1'b0,  10'd19},{  8'd0, 1'b0,  10'd34},{  8'd0, 1'b0,  10'd44},{  8'd0, 1'b0,  10'd49},{  8'd0, 1'b0,  10'd54},{  8'd0, 1'b0,  10'd59},{  8'd0, 1'b0, 10'd109},{  8'd0, 1'b0, 10'd114},{  8'd0, 1'b0, 10'd124},{  8'd0, 1'b0, 10'd129},{  8'd0, 1'b1, 10'd144}
};
localparam int          cSHORT_HS_TAB_7BY15_PACKED_SIZE = 203;
localparam bit [18 : 0] cSHORT_HS_TAB_7BY15_PACKED[cSHORT_HS_TAB_7BY15_PACKED_SIZE] = '{
{  1'b0, 1'b0,  8'd22,    9'd0},{  1'b0, 1'b0,  8'd21,    9'd0},{  1'b0, 1'b0,  8'd18,  9'd302},{  1'b0, 1'b0,   8'd7,  9'd327},{  1'b0, 1'b0,   8'd3,  9'd113},{  1'b0, 1'b0,   8'd2,   9'd59},{  1'b0, 1'b0,   8'd1,  9'd251},{  1'b0, 1'b1,   8'd0,  9'd134},
{  1'b0, 1'b0,  8'd23,    9'd0},{  1'b0, 1'b0,  8'd22,    9'd0},{  1'b0, 1'b0,  8'd13,  9'd220},{  1'b0, 1'b0,  8'd10,  9'd358},{  1'b0, 1'b0,   8'd3,  9'd262},{  1'b0, 1'b0,   8'd2,  9'd355},{  1'b0, 1'b0,   8'd1,  9'd335},{  1'b0, 1'b1,   8'd0,   9'd13},
{  1'b0, 1'b0,  8'd24,    9'd0},{  1'b0, 1'b0,  8'd23,    9'd0},{  1'b0, 1'b0,  8'd16,  9'd345},{  1'b0, 1'b0,  8'd10,  9'd108},{  1'b0, 1'b0,   8'd3,  9'd144},{  1'b0, 1'b0,   8'd2,  9'd201},{  1'b0, 1'b0,   8'd1,  9'd258},{  1'b0, 1'b1,   8'd0,    9'd0},
{  1'b0, 1'b0,  8'd26,    9'd0},{  1'b0, 1'b0,  8'd25,    9'd0},{  1'b0, 1'b0,  8'd16,    9'd8},{  1'b0, 1'b0,  8'd11,  9'd314},{  1'b0, 1'b0,   8'd3,  9'd240},{  1'b0, 1'b0,   8'd2,  9'd336},{  1'b0, 1'b0,   8'd1,  9'd179},{  1'b0, 1'b1,   8'd0,  9'd171},
{  1'b0, 1'b0,  8'd27,    9'd0},{  1'b0, 1'b0,  8'd26,    9'd0},{  1'b0, 1'b0,  8'd18,  9'd314},{  1'b0, 1'b0,  8'd10,  9'd310},{  1'b0, 1'b0,   8'd3,  9'd345},{  1'b0, 1'b0,   8'd2,  9'd338},{  1'b0, 1'b0,   8'd1,  9'd349},{  1'b0, 1'b1,   8'd0,  9'd355},
{  1'b0, 1'b0,  8'd33,    9'd0},{  1'b0, 1'b0,  8'd32,    9'd0},{  1'b0, 1'b0,  8'd19,   9'd89},{  1'b0, 1'b0,   8'd7,   9'd92},{  1'b0, 1'b0,   8'd3,  9'd123},{  1'b0, 1'b0,   8'd2,  9'd313},{  1'b0, 1'b0,   8'd1,  9'd263},{  1'b0, 1'b1,   8'd0,   9'd84},
{  1'b0, 1'b0,  8'd34,    9'd0},{  1'b0, 1'b0,  8'd33,    9'd0},{  1'b0, 1'b0,  8'd20,  9'd208},{  1'b0, 1'b0,  8'd11,   9'd87},{  1'b0, 1'b0,   8'd3,  9'd231},{  1'b0, 1'b0,   8'd2,  9'd158},{  1'b0, 1'b0,   8'd1,  9'd284},{  1'b0, 1'b1,   8'd0,   9'd66},
{  1'b0, 1'b0,  8'd35,    9'd0},{  1'b0, 1'b0,  8'd34,    9'd0},{  1'b0, 1'b0,  8'd14,  9'd349},{  1'b0, 1'b0,   8'd6,  9'd170},{  1'b0, 1'b0,   8'd3,  9'd113},{  1'b0, 1'b0,   8'd2,  9'd357},{  1'b0, 1'b0,   8'd1,  9'd278},{  1'b0, 1'b1,   8'd0,  9'd324},
{  1'b0, 1'b0,  8'd37,    9'd0},{  1'b0, 1'b0,  8'd36,    9'd0},{  1'b0, 1'b0,  8'd20,   9'd40},{  1'b0, 1'b0,   8'd8,  9'd290},{  1'b0, 1'b0,   8'd3,  9'd285},{  1'b0, 1'b0,   8'd2,  9'd248},{  1'b0, 1'b0,   8'd1,  9'd128},{  1'b0, 1'b1,   8'd0,  9'd308},
{  1'b0, 1'b0,  8'd39,    9'd0},{  1'b0, 1'b0,  8'd38,    9'd0},{  1'b0, 1'b0,  8'd18,   9'd37},{  1'b0, 1'b0,  8'd11,  9'd154},{  1'b0, 1'b0,   8'd3,   9'd29},{  1'b0, 1'b0,   8'd2,    9'd0},{  1'b0, 1'b0,   8'd1,  9'd265},{  1'b0, 1'b1,   8'd0,  9'd297},
{  1'b0, 1'b0,  8'd40,    9'd0},{  1'b0, 1'b0,  8'd39,    9'd0},{  1'b0, 1'b0,  8'd14,  9'd244},{  1'b0, 1'b0,   8'd9,  9'd324},{  1'b0, 1'b0,   8'd3,  9'd355},{  1'b0, 1'b0,   8'd2,    9'd7},{  1'b0, 1'b0,   8'd1,  9'd357},{  1'b0, 1'b1,   8'd0,  9'd126},
{  1'b0, 1'b0,  8'd42,    9'd0},{  1'b0, 1'b0,  8'd41,    9'd0},{  1'b0, 1'b0,  8'd16,  9'd193},{  1'b0, 1'b0,  8'd10,   9'd58},{  1'b0, 1'b0,   8'd3,  9'd273},{  1'b0, 1'b0,   8'd2,  9'd194},{  1'b0, 1'b0,   8'd1,   9'd49},{  1'b0, 1'b1,   8'd0,  9'd328},
{  1'b0, 1'b0,  8'd43,    9'd0},{  1'b0, 1'b0,  8'd42,    9'd0},{  1'b0, 1'b0,  8'd17,   9'd24},{  1'b0, 1'b0,   8'd8,   9'd41},{  1'b0, 1'b0,   8'd3,  9'd138},{  1'b0, 1'b0,   8'd2,  9'd145},{  1'b0, 1'b0,   8'd1,  9'd314},{  1'b0, 1'b1,   8'd0,  9'd359},
{  1'b1, 1'b0,  8'd44,    9'd1},{  1'b0, 1'b0,  8'd21,    9'd0},{  1'b0, 1'b0,  8'd13,  9'd131},{  1'b0, 1'b0,   8'd9,  9'd252},{  1'b0, 1'b0,   8'd5,  9'd125},{  1'b0, 1'b0,   8'd3,  9'd352},{  1'b0, 1'b0,   8'd2,   9'd97},{  1'b0, 1'b0,   8'd1,  9'd113},{  1'b0, 1'b1,   8'd0,  9'd359},
{  1'b0, 1'b0,  8'd25,    9'd0},{  1'b0, 1'b0,  8'd24,    9'd0},{  1'b0, 1'b0,  8'd13,  9'd193},{  1'b0, 1'b0,   8'd7,  9'd356},{  1'b0, 1'b0,   8'd4,  9'd337},{  1'b0, 1'b0,   8'd3,  9'd134},{  1'b0, 1'b0,   8'd2,  9'd267},{  1'b0, 1'b0,   8'd1,  9'd211},{  1'b0, 1'b1,   8'd0,  9'd299},
{  1'b0, 1'b0,  8'd28,    9'd0},{  1'b0, 1'b0,  8'd27,    9'd0},{  1'b0, 1'b0,  8'd15,  9'd332},{  1'b0, 1'b0,   8'd8,  9'd135},{  1'b0, 1'b0,   8'd4,  9'd359},{  1'b0, 1'b0,   8'd3,  9'd127},{  1'b0, 1'b0,   8'd2,  9'd231},{  1'b0, 1'b0,   8'd1,   9'd79},{  1'b0, 1'b1,   8'd0,  9'd272},
{  1'b0, 1'b0,  8'd29,    9'd0},{  1'b0, 1'b0,  8'd28,    9'd0},{  1'b0, 1'b0,  8'd17,  9'd359},{  1'b0, 1'b0,   8'd8,  9'd107},{  1'b0, 1'b0,   8'd5,    9'd2},{  1'b0, 1'b0,   8'd3,  9'd349},{  1'b0, 1'b0,   8'd2,  9'd332},{  1'b0, 1'b0,   8'd1,   9'd50},{  1'b0, 1'b1,   8'd0,  9'd273},
{  1'b0, 1'b0,  8'd30,    9'd0},{  1'b0, 1'b0,  8'd29,    9'd0},{  1'b0, 1'b0,  8'd20,   9'd83},{  1'b0, 1'b0,  8'd12,  9'd248},{  1'b0, 1'b0,   8'd6,   9'd75},{  1'b0, 1'b0,   8'd3,  9'd243},{  1'b0, 1'b0,   8'd2,  9'd281},{  1'b0, 1'b0,   8'd1,  9'd147},{  1'b0, 1'b1,   8'd0,  9'd346},
{  1'b0, 1'b0,  8'd31,    9'd0},{  1'b0, 1'b0,  8'd30,    9'd0},{  1'b0, 1'b0,  8'd15,  9'd138},{  1'b0, 1'b0,  8'd12,    9'd0},{  1'b0, 1'b0,   8'd5,  9'd343},{  1'b0, 1'b0,   8'd3,  9'd324},{  1'b0, 1'b0,   8'd2,  9'd266},{  1'b0, 1'b0,   8'd1,  9'd358},{  1'b0, 1'b1,   8'd0,  9'd257},
{  1'b0, 1'b0,  8'd32,    9'd0},{  1'b0, 1'b0,  8'd31,    9'd0},{  1'b0, 1'b0,  8'd19,  9'd341},{  1'b0, 1'b0,  8'd11,  9'd355},{  1'b0, 1'b0,   8'd5,   9'd81},{  1'b0, 1'b0,   8'd3,  9'd267},{  1'b0, 1'b0,   8'd2,   9'd46},{  1'b0, 1'b0,   8'd1,  9'd170},{  1'b0, 1'b1,   8'd0,  9'd338},
{  1'b0, 1'b0,  8'd36,    9'd0},{  1'b0, 1'b0,  8'd35,    9'd0},{  1'b0, 1'b0,  8'd15,  9'd217},{  1'b0, 1'b0,   8'd9,  9'd345},{  1'b0, 1'b0,   8'd4,  9'd330},{  1'b0, 1'b0,   8'd3,  9'd356},{  1'b0, 1'b0,   8'd2,  9'd320},{  1'b0, 1'b0,   8'd1,   9'd76},{  1'b0, 1'b1,   8'd0,   9'd13},
{  1'b0, 1'b0,  8'd38,    9'd0},{  1'b0, 1'b0,  8'd37,    9'd0},{  1'b0, 1'b0,  8'd17,  9'd224},{  1'b0, 1'b0,   8'd9,   9'd90},{  1'b0, 1'b0,   8'd6,  9'd353},{  1'b0, 1'b0,   8'd3,  9'd330},{  1'b0, 1'b0,   8'd2,  9'd298},{  1'b0, 1'b0,   8'd1,  9'd322},{  1'b0, 1'b1,   8'd0,    9'd5},
{  1'b0, 1'b0,  8'd41,    9'd0},{  1'b0, 1'b0,  8'd40,    9'd0},{  1'b0, 1'b0,  8'd14,  9'd237},{  1'b0, 1'b0,  8'd12,  9'd311},{  1'b0, 1'b0,   8'd4,  9'd143},{  1'b0, 1'b0,   8'd3,  9'd339},{  1'b0, 1'b0,   8'd2,   9'd95},{  1'b0, 1'b0,   8'd1,   9'd14},{  1'b0, 1'b1,   8'd0,  9'd250},
{  1'b0, 1'b0,  8'd44,    9'd0},{  1'b0, 1'b0,  8'd43,    9'd0},{  1'b0, 1'b0,  8'd19,   9'd50},{  1'b0, 1'b0,   8'd7,  9'd268},{  1'b0, 1'b0,   8'd6,  9'd332},{  1'b0, 1'b0,   8'd3,  9'd346},{  1'b0, 1'b0,   8'd2,   9'd60},{  1'b0, 1'b0,   8'd1,  9'd204},{  1'b0, 1'b1,   8'd0,   9'd40}
};
localparam bit [18 : 0] cSHORT_HS_V_TAB_7BY15_PACKED[cSHORT_HS_TAB_7BY15_PACKED_SIZE] = '{
{ 8'd44, 1'b0, 10'd104},{ 8'd44, 1'b1, 10'd194},
{ 8'd43, 1'b0,  10'd96},{ 8'd43, 1'b1, 10'd195},
{ 8'd42, 1'b0,  10'd88},{ 8'd42, 1'b1,  10'd97},
{ 8'd41, 1'b0, 10'd185},{ 8'd41, 1'b1,  10'd89},
{ 8'd40, 1'b0,  10'd80},{ 8'd40, 1'b1, 10'd186},
{ 8'd39, 1'b0,  10'd72},{ 8'd39, 1'b1,  10'd81},
{ 8'd38, 1'b0, 10'd176},{ 8'd38, 1'b1,  10'd73},
{ 8'd37, 1'b0,  10'd64},{ 8'd37, 1'b1, 10'd177},
{ 8'd36, 1'b0, 10'd167},{ 8'd36, 1'b1,  10'd65},
{ 8'd35, 1'b0,  10'd56},{ 8'd35, 1'b1, 10'd168},
{ 8'd34, 1'b0,  10'd48},{ 8'd34, 1'b1,  10'd57},
{ 8'd33, 1'b0,  10'd40},{ 8'd33, 1'b1,  10'd49},
{ 8'd32, 1'b0, 10'd158},{ 8'd32, 1'b1,  10'd41},
{ 8'd31, 1'b0, 10'd149},{ 8'd31, 1'b1, 10'd159},
{ 8'd30, 1'b0, 10'd140},{ 8'd30, 1'b1, 10'd150},
{ 8'd29, 1'b0, 10'd131},{ 8'd29, 1'b1, 10'd141},
{ 8'd28, 1'b0, 10'd122},{ 8'd28, 1'b1, 10'd132},
{ 8'd27, 1'b0,  10'd32},{ 8'd27, 1'b1, 10'd123},
{ 8'd26, 1'b0,  10'd24},{ 8'd26, 1'b1,  10'd33},
{ 8'd25, 1'b0, 10'd113},{ 8'd25, 1'b1,  10'd25},
{ 8'd24, 1'b0,  10'd16},{ 8'd24, 1'b1, 10'd114},
{ 8'd23, 1'b0,   10'd8},{ 8'd23, 1'b1,  10'd17},
{ 8'd22, 1'b0,   10'd0},{ 8'd22, 1'b1,   10'd9},
{ 8'd21, 1'b0, 10'd105},{ 8'd21, 1'b1,   10'd1},
{ 8'd20, 1'b0, 10'd142},{ 8'd20, 1'b0,  10'd50},{ 8'd20, 1'b1,  10'd66},
{ 8'd19, 1'b0, 10'd160},{ 8'd19, 1'b0,  10'd42},{ 8'd19, 1'b1, 10'd196},
{ 8'd18, 1'b0,   10'd2},{ 8'd18, 1'b0,  10'd34},{ 8'd18, 1'b1,  10'd74},
{ 8'd17, 1'b0, 10'd133},{ 8'd17, 1'b0, 10'd178},{ 8'd17, 1'b1,  10'd98},
{ 8'd16, 1'b0,  10'd18},{ 8'd16, 1'b0,  10'd26},{ 8'd16, 1'b1,  10'd90},
{ 8'd15, 1'b0, 10'd124},{ 8'd15, 1'b0, 10'd151},{ 8'd15, 1'b1, 10'd169},
{ 8'd14, 1'b0,  10'd58},{ 8'd14, 1'b0,  10'd82},{ 8'd14, 1'b1, 10'd187},
{ 8'd13, 1'b0, 10'd106},{ 8'd13, 1'b0,  10'd10},{ 8'd13, 1'b1, 10'd115},
{ 8'd12, 1'b0, 10'd143},{ 8'd12, 1'b0, 10'd152},{ 8'd12, 1'b1, 10'd188},
{ 8'd11, 1'b0,  10'd27},{ 8'd11, 1'b0, 10'd161},{ 8'd11, 1'b0,  10'd51},{ 8'd11, 1'b1,  10'd75},
{ 8'd10, 1'b0,  10'd11},{ 8'd10, 1'b0,  10'd19},{ 8'd10, 1'b0,  10'd35},{ 8'd10, 1'b1,  10'd91},
{  8'd9, 1'b0, 10'd107},{  8'd9, 1'b0, 10'd170},{  8'd9, 1'b0, 10'd179},{  8'd9, 1'b1,  10'd83},
{  8'd8, 1'b0, 10'd125},{  8'd8, 1'b0, 10'd134},{  8'd8, 1'b0,  10'd67},{  8'd8, 1'b1,  10'd99},
{  8'd7, 1'b0,   10'd3},{  8'd7, 1'b0, 10'd116},{  8'd7, 1'b0,  10'd43},{  8'd7, 1'b1, 10'd197},
{  8'd6, 1'b0, 10'd144},{  8'd6, 1'b0,  10'd59},{  8'd6, 1'b0, 10'd180},{  8'd6, 1'b1, 10'd198},
{  8'd5, 1'b0, 10'd108},{  8'd5, 1'b0, 10'd135},{  8'd5, 1'b0, 10'd153},{  8'd5, 1'b1, 10'd162},
{  8'd4, 1'b0, 10'd117},{  8'd4, 1'b0, 10'd126},{  8'd4, 1'b0, 10'd171},{  8'd4, 1'b1, 10'd189},
{  8'd3, 1'b0, 10'd109},{  8'd3, 1'b0,   10'd4},{  8'd3, 1'b0,  10'd12},{  8'd3, 1'b0,  10'd20},{  8'd3, 1'b0, 10'd118},{  8'd3, 1'b0,  10'd28},{  8'd3, 1'b0,  10'd36},{  8'd3, 1'b0, 10'd127},{  8'd3, 1'b0, 10'd136},{  8'd3, 1'b0, 10'd145},{  8'd3, 1'b0, 10'd154},{  8'd3, 1'b0, 10'd163},{  8'd3, 1'b0,  10'd44},{  8'd3, 1'b0,  10'd52},{  8'd3, 1'b0,  10'd60},{  8'd3, 1'b0, 10'd172},{  8'd3, 1'b0,  10'd68},{  8'd3, 1'b0, 10'd181},{  8'd3, 1'b0,  10'd76},{  8'd3, 1'b0,  10'd84},{  8'd3, 1'b0, 10'd190},{  8'd3, 1'b0,  10'd92},{  8'd3, 1'b0, 10'd100},{  8'd3, 1'b1, 10'd199},
{  8'd2, 1'b0, 10'd110},{  8'd2, 1'b0,   10'd5},{  8'd2, 1'b0,  10'd13},{  8'd2, 1'b0,  10'd21},{  8'd2, 1'b0, 10'd119},{  8'd2, 1'b0,  10'd29},{  8'd2, 1'b0,  10'd37},{  8'd2, 1'b0, 10'd128},{  8'd2, 1'b0, 10'd137},{  8'd2, 1'b0, 10'd146},{  8'd2, 1'b0, 10'd155},{  8'd2, 1'b0, 10'd164},{  8'd2, 1'b0,  10'd45},{  8'd2, 1'b0,  10'd53},{  8'd2, 1'b0,  10'd61},{  8'd2, 1'b0, 10'd173},{  8'd2, 1'b0,  10'd69},{  8'd2, 1'b0, 10'd182},{  8'd2, 1'b0,  10'd77},{  8'd2, 1'b0,  10'd85},{  8'd2, 1'b0, 10'd191},{  8'd2, 1'b0,  10'd93},{  8'd2, 1'b0, 10'd101},{  8'd2, 1'b1, 10'd200},
{  8'd1, 1'b0, 10'd111},{  8'd1, 1'b0,   10'd6},{  8'd1, 1'b0,  10'd14},{  8'd1, 1'b0,  10'd22},{  8'd1, 1'b0, 10'd120},{  8'd1, 1'b0,  10'd30},{  8'd1, 1'b0,  10'd38},{  8'd1, 1'b0, 10'd129},{  8'd1, 1'b0, 10'd138},{  8'd1, 1'b0, 10'd147},{  8'd1, 1'b0, 10'd156},{  8'd1, 1'b0, 10'd165},{  8'd1, 1'b0,  10'd46},{  8'd1, 1'b0,  10'd54},{  8'd1, 1'b0,  10'd62},{  8'd1, 1'b0, 10'd174},{  8'd1, 1'b0,  10'd70},{  8'd1, 1'b0, 10'd183},{  8'd1, 1'b0,  10'd78},{  8'd1, 1'b0,  10'd86},{  8'd1, 1'b0, 10'd192},{  8'd1, 1'b0,  10'd94},{  8'd1, 1'b0, 10'd102},{  8'd1, 1'b1, 10'd201},
{  8'd0, 1'b0, 10'd112},{  8'd0, 1'b0,   10'd7},{  8'd0, 1'b0,  10'd15},{  8'd0, 1'b0,  10'd23},{  8'd0, 1'b0, 10'd121},{  8'd0, 1'b0,  10'd31},{  8'd0, 1'b0,  10'd39},{  8'd0, 1'b0, 10'd130},{  8'd0, 1'b0, 10'd139},{  8'd0, 1'b0, 10'd148},{  8'd0, 1'b0, 10'd157},{  8'd0, 1'b0, 10'd166},{  8'd0, 1'b0,  10'd47},{  8'd0, 1'b0,  10'd55},{  8'd0, 1'b0,  10'd63},{  8'd0, 1'b0, 10'd175},{  8'd0, 1'b0,  10'd71},{  8'd0, 1'b0, 10'd184},{  8'd0, 1'b0,  10'd79},{  8'd0, 1'b0,  10'd87},{  8'd0, 1'b0, 10'd193},{  8'd0, 1'b0,  10'd95},{  8'd0, 1'b0, 10'd103},{  8'd0, 1'b1, 10'd202}
};
localparam int          cSHORT_HS_TAB_8BY15_PACKED_SIZE = 209;
localparam bit [18 : 0] cSHORT_HS_TAB_8BY15_PACKED[cSHORT_HS_TAB_8BY15_PACKED_SIZE] = '{
{  1'b0, 1'b0,  8'd41,    9'd0},{  1'b0, 1'b0,  8'd40,    9'd0},{  1'b0, 1'b0,  8'd20,  9'd103},{  1'b0, 1'b0,  8'd16,  9'd280},{  1'b0, 1'b0,   8'd4,  9'd308},{  1'b0, 1'b0,   8'd3,  9'd277},{  1'b0, 1'b0,   8'd2,  9'd199},{  1'b0, 1'b0,   8'd1,  9'd236},{  1'b0, 1'b1,   8'd0,  9'd338},
{  1'b1, 1'b0,  8'd44,    9'd1},{  1'b0, 1'b0,  8'd24,    9'd0},{  1'b0, 1'b0,  8'd21,  9'd101},{  1'b0, 1'b0,  8'd13,  9'd349},{  1'b0, 1'b0,   8'd6,  9'd245},{  1'b0, 1'b0,   8'd4,  9'd138},{  1'b0, 1'b0,   8'd3,  9'd322},{  1'b0, 1'b0,   8'd2,  9'd343},{  1'b0, 1'b0,   8'd1,  9'd356},{  1'b0, 1'b1,   8'd0,  9'd222},
{  1'b0, 1'b0,  8'd25,    9'd0},{  1'b0, 1'b0,  8'd24,    9'd0},{  1'b0, 1'b0,  8'd22,  9'd148},{  1'b0, 1'b0,  8'd14,  9'd132},{  1'b0, 1'b0,   8'd5,  9'd194},{  1'b0, 1'b0,   8'd4,  9'd219},{  1'b0, 1'b0,   8'd3,  9'd133},{  1'b0, 1'b0,   8'd2,  9'd277},{  1'b0, 1'b0,   8'd1,  9'd333},{  1'b0, 1'b1,   8'd0,  9'd238},
{  1'b0, 1'b0,  8'd26,    9'd0},{  1'b0, 1'b0,  8'd25,    9'd0},{  1'b0, 1'b0,  8'd19,  9'd353},{  1'b0, 1'b0,  8'd12,  9'd272},{  1'b0, 1'b0,   8'd8,  9'd244},{  1'b0, 1'b0,   8'd4,  9'd355},{  1'b0, 1'b0,   8'd3,  9'd281},{  1'b0, 1'b0,   8'd2,  9'd287},{  1'b0, 1'b0,   8'd1,  9'd338},{  1'b0, 1'b1,   8'd0,   9'd94},
{  1'b0, 1'b0,  8'd27,    9'd0},{  1'b0, 1'b0,  8'd26,    9'd0},{  1'b0, 1'b0,  8'd19,  9'd326},{  1'b0, 1'b0,  8'd11,  9'd257},{  1'b0, 1'b0,   8'd9,  9'd290},{  1'b0, 1'b0,   8'd4,   9'd32},{  1'b0, 1'b0,   8'd3,  9'd323},{  1'b0, 1'b0,   8'd2,  9'd279},{  1'b0, 1'b0,   8'd1,   9'd85},{  1'b0, 1'b1,   8'd0,   9'd28},
{  1'b0, 1'b0,  8'd28,    9'd0},{  1'b0, 1'b0,  8'd27,    9'd0},{  1'b0, 1'b0,  8'd20,  9'd359},{  1'b0, 1'b0,  8'd15,  9'd140},{  1'b0, 1'b0,   8'd9,  9'd135},{  1'b0, 1'b0,   8'd4,   9'd39},{  1'b0, 1'b0,   8'd3,  9'd316},{  1'b0, 1'b0,   8'd2,  9'd257},{  1'b0, 1'b0,   8'd1,  9'd356},{  1'b0, 1'b1,   8'd0,   9'd95},
{  1'b0, 1'b0,  8'd29,    9'd0},{  1'b0, 1'b0,  8'd28,    9'd0},{  1'b0, 1'b0,  8'd19,   9'd76},{  1'b0, 1'b0,  8'd16,  9'd220},{  1'b0, 1'b0,   8'd5,  9'd348},{  1'b0, 1'b0,   8'd4,  9'd343},{  1'b0, 1'b0,   8'd3,  9'd353},{  1'b0, 1'b0,   8'd2,  9'd284},{  1'b0, 1'b0,   8'd1,  9'd328},{  1'b0, 1'b1,   8'd0,  9'd173},
{  1'b0, 1'b0,  8'd30,    9'd0},{  1'b0, 1'b0,  8'd29,    9'd0},{  1'b0, 1'b0,  8'd22,  9'd240},{  1'b0, 1'b0,  8'd12,  9'd246},{  1'b0, 1'b0,   8'd7,  9'd152},{  1'b0, 1'b0,   8'd4,   9'd44},{  1'b0, 1'b0,   8'd3,  9'd160},{  1'b0, 1'b0,   8'd2,  9'd255},{  1'b0, 1'b0,   8'd1,  9'd272},{  1'b0, 1'b1,   8'd0,   9'd18},
{  1'b0, 1'b0,  8'd31,    9'd0},{  1'b0, 1'b0,  8'd30,    9'd0},{  1'b0, 1'b0,  8'd23,   9'd48},{  1'b0, 1'b0,  8'd15,  9'd128},{  1'b0, 1'b0,   8'd7,  9'd231},{  1'b0, 1'b0,   8'd4,  9'd355},{  1'b0, 1'b0,   8'd3,   9'd27},{  1'b0, 1'b0,   8'd2,  9'd297},{  1'b0, 1'b0,   8'd1,  9'd352},{  1'b0, 1'b1,   8'd0,  9'd342},
{  1'b0, 1'b0,  8'd32,    9'd0},{  1'b0, 1'b0,  8'd31,    9'd0},{  1'b0, 1'b0,  8'd18,  9'd350},{  1'b0, 1'b0,  8'd16,  9'd153},{  1'b0, 1'b0,   8'd6,  9'd340},{  1'b0, 1'b0,   8'd4,   9'd42},{  1'b0, 1'b0,   8'd3,  9'd335},{  1'b0, 1'b0,   8'd2,  9'd139},{  1'b0, 1'b0,   8'd1,  9'd278},{  1'b0, 1'b1,   8'd0,  9'd246},
{  1'b0, 1'b0,  8'd33,    9'd0},{  1'b0, 1'b0,  8'd32,    9'd0},{  1'b0, 1'b0,  8'd23,  9'd355},{  1'b0, 1'b0,  8'd12,   9'd98},{  1'b0, 1'b0,   8'd5,  9'd199},{  1'b0, 1'b0,   8'd4,   9'd62},{  1'b0, 1'b0,   8'd3,  9'd277},{  1'b0, 1'b0,   8'd2,  9'd316},{  1'b0, 1'b0,   8'd1,  9'd267},{  1'b0, 1'b1,   8'd0,  9'd271},
{  1'b0, 1'b0,  8'd34,    9'd0},{  1'b0, 1'b0,  8'd33,    9'd0},{  1'b0, 1'b0,  8'd17,   9'd80},{  1'b0, 1'b0,  8'd14,   9'd85},{  1'b0, 1'b0,   8'd6,  9'd357},{  1'b0, 1'b0,   8'd4,    9'd8},{  1'b0, 1'b0,   8'd3,  9'd159},{  1'b0, 1'b0,   8'd2,  9'd134},{  1'b0, 1'b0,   8'd1,  9'd214},{  1'b0, 1'b1,   8'd0,   9'd20},
{  1'b0, 1'b0,  8'd35,    9'd0},{  1'b0, 1'b0,  8'd34,    9'd0},{  1'b0, 1'b0,  8'd17,  9'd291},{  1'b0, 1'b0,  8'd10,    9'd0},{  1'b0, 1'b0,   8'd7,  9'd332},{  1'b0, 1'b0,   8'd4,  9'd347},{  1'b0, 1'b0,   8'd3,   9'd98},{  1'b0, 1'b0,   8'd2,  9'd331},{  1'b0, 1'b0,   8'd1,  9'd346},{  1'b0, 1'b1,   8'd0,    9'd1},
{  1'b0, 1'b0,  8'd36,    9'd0},{  1'b0, 1'b0,  8'd35,    9'd0},{  1'b0, 1'b0,  8'd17,  9'd324},{  1'b0, 1'b0,  8'd13,  9'd341},{  1'b0, 1'b0,   8'd6,  9'd286},{  1'b0, 1'b0,   8'd4,   9'd57},{  1'b0, 1'b0,   8'd3,   9'd69},{  1'b0, 1'b0,   8'd2,  9'd228},{  1'b0, 1'b0,   8'd1,   9'd89},{  1'b0, 1'b1,   8'd0,  9'd103},
{  1'b0, 1'b0,  8'd37,    9'd0},{  1'b0, 1'b0,  8'd36,    9'd0},{  1'b0, 1'b0,  8'd21,  9'd325},{  1'b0, 1'b0,  8'd14,  9'd166},{  1'b0, 1'b0,   8'd8,  9'd328},{  1'b0, 1'b0,   8'd4,  9'd206},{  1'b0, 1'b0,   8'd3,  9'd326},{  1'b0, 1'b0,   8'd2,  9'd235},{  1'b0, 1'b0,   8'd1,  9'd310},{  1'b0, 1'b1,   8'd0,  9'd213},
{  1'b0, 1'b0,  8'd38,    9'd0},{  1'b0, 1'b0,  8'd37,    9'd0},{  1'b0, 1'b0,  8'd18,  9'd325},{  1'b0, 1'b0,  8'd11,  9'd344},{  1'b0, 1'b0,   8'd5,  9'd359},{  1'b0, 1'b0,   8'd4,    9'd0},{  1'b0, 1'b0,   8'd3,  9'd113},{  1'b0, 1'b0,   8'd2,  9'd204},{  1'b0, 1'b0,   8'd1,  9'd234},{  1'b0, 1'b1,   8'd0,  9'd200},
{  1'b0, 1'b0,  8'd39,    9'd0},{  1'b0, 1'b0,  8'd38,    9'd0},{  1'b0, 1'b0,  8'd18,  9'd238},{  1'b0, 1'b0,  8'd15,  9'd320},{  1'b0, 1'b0,   8'd9,  9'd336},{  1'b0, 1'b0,   8'd4,  9'd343},{  1'b0, 1'b0,   8'd3,  9'd359},{  1'b0, 1'b0,   8'd2,  9'd347},{  1'b0, 1'b0,   8'd1,  9'd129},{  1'b0, 1'b1,   8'd0,   9'd61},
{  1'b0, 1'b0,  8'd40,    9'd0},{  1'b0, 1'b0,  8'd39,    9'd0},{  1'b0, 1'b0,  8'd22,   9'd92},{  1'b0, 1'b0,  8'd10,  9'd257},{  1'b0, 1'b0,   8'd9,  9'd354},{  1'b0, 1'b0,   8'd4,  9'd247},{  1'b0, 1'b0,   8'd3,  9'd235},{  1'b0, 1'b0,   8'd2,  9'd358},{  1'b0, 1'b0,   8'd1,  9'd270},{  1'b0, 1'b1,   8'd0,  9'd101},
{  1'b0, 1'b0,  8'd42,    9'd0},{  1'b0, 1'b0,  8'd41,    9'd0},{  1'b0, 1'b0,  8'd20,  9'd351},{  1'b0, 1'b0,  8'd10,  9'd177},{  1'b0, 1'b0,   8'd8,  9'd267},{  1'b0, 1'b0,   8'd4,  9'd311},{  1'b0, 1'b0,   8'd3,  9'd353},{  1'b0, 1'b0,   8'd2,  9'd270},{  1'b0, 1'b0,   8'd1,  9'd336},{  1'b0, 1'b1,   8'd0,  9'd331},
{  1'b0, 1'b0,  8'd43,    9'd0},{  1'b0, 1'b0,  8'd42,    9'd0},{  1'b0, 1'b0,  8'd21,  9'd335},{  1'b0, 1'b0,  8'd11,  9'd118},{  1'b0, 1'b0,   8'd7,  9'd334},{  1'b0, 1'b0,   8'd4,  9'd331},{  1'b0, 1'b0,   8'd3,   9'd97},{  1'b0, 1'b0,   8'd2,  9'd132},{  1'b0, 1'b0,   8'd1,  9'd358},{  1'b0, 1'b1,   8'd0,  9'd339},
{  1'b0, 1'b0,  8'd44,    9'd0},{  1'b0, 1'b0,  8'd43,    9'd0},{  1'b0, 1'b0,  8'd23,   9'd12},{  1'b0, 1'b0,  8'd13,   9'd89},{  1'b0, 1'b0,   8'd8,  9'd150},{  1'b0, 1'b0,   8'd4,  9'd354},{  1'b0, 1'b0,   8'd3,   9'd86},{  1'b0, 1'b0,   8'd2,  9'd354},{  1'b0, 1'b0,   8'd1,   9'd90},{  1'b0, 1'b1,   8'd0,  9'd204}
};
localparam bit [18 : 0] cSHORT_HS_V_TAB_8BY15_PACKED[cSHORT_HS_TAB_8BY15_PACKED_SIZE] = '{
{ 8'd44, 1'b0,   10'd9},{ 8'd44, 1'b1, 10'd199},
{ 8'd43, 1'b0, 10'd189},{ 8'd43, 1'b1, 10'd200},
{ 8'd42, 1'b0, 10'd179},{ 8'd42, 1'b1, 10'd190},
{ 8'd41, 1'b0,   10'd0},{ 8'd41, 1'b1, 10'd180},
{ 8'd40, 1'b0, 10'd169},{ 8'd40, 1'b1,   10'd1},
{ 8'd39, 1'b0, 10'd159},{ 8'd39, 1'b1, 10'd170},
{ 8'd38, 1'b0, 10'd149},{ 8'd38, 1'b1, 10'd160},
{ 8'd37, 1'b0, 10'd139},{ 8'd37, 1'b1, 10'd150},
{ 8'd36, 1'b0, 10'd129},{ 8'd36, 1'b1, 10'd140},
{ 8'd35, 1'b0, 10'd119},{ 8'd35, 1'b1, 10'd130},
{ 8'd34, 1'b0, 10'd109},{ 8'd34, 1'b1, 10'd120},
{ 8'd33, 1'b0,  10'd99},{ 8'd33, 1'b1, 10'd110},
{ 8'd32, 1'b0,  10'd89},{ 8'd32, 1'b1, 10'd100},
{ 8'd31, 1'b0,  10'd79},{ 8'd31, 1'b1,  10'd90},
{ 8'd30, 1'b0,  10'd69},{ 8'd30, 1'b1,  10'd80},
{ 8'd29, 1'b0,  10'd59},{ 8'd29, 1'b1,  10'd70},
{ 8'd28, 1'b0,  10'd49},{ 8'd28, 1'b1,  10'd60},
{ 8'd27, 1'b0,  10'd39},{ 8'd27, 1'b1,  10'd50},
{ 8'd26, 1'b0,  10'd29},{ 8'd26, 1'b1,  10'd40},
{ 8'd25, 1'b0,  10'd19},{ 8'd25, 1'b1,  10'd30},
{ 8'd24, 1'b0,  10'd10},{ 8'd24, 1'b1,  10'd20},
{ 8'd23, 1'b0,  10'd81},{ 8'd23, 1'b0, 10'd101},{ 8'd23, 1'b1, 10'd201},
{ 8'd22, 1'b0,  10'd21},{ 8'd22, 1'b0,  10'd71},{ 8'd22, 1'b1, 10'd171},
{ 8'd21, 1'b0,  10'd11},{ 8'd21, 1'b0, 10'd141},{ 8'd21, 1'b1, 10'd191},
{ 8'd20, 1'b0,  10'd51},{ 8'd20, 1'b0,   10'd2},{ 8'd20, 1'b1, 10'd181},
{ 8'd19, 1'b0,  10'd31},{ 8'd19, 1'b0,  10'd41},{ 8'd19, 1'b1,  10'd61},
{ 8'd18, 1'b0,  10'd91},{ 8'd18, 1'b0, 10'd151},{ 8'd18, 1'b1, 10'd161},
{ 8'd17, 1'b0, 10'd111},{ 8'd17, 1'b0, 10'd121},{ 8'd17, 1'b1, 10'd131},
{ 8'd16, 1'b0,  10'd62},{ 8'd16, 1'b0,  10'd92},{ 8'd16, 1'b1,   10'd3},
{ 8'd15, 1'b0,  10'd52},{ 8'd15, 1'b0,  10'd82},{ 8'd15, 1'b1, 10'd162},
{ 8'd14, 1'b0,  10'd22},{ 8'd14, 1'b0, 10'd112},{ 8'd14, 1'b1, 10'd142},
{ 8'd13, 1'b0,  10'd12},{ 8'd13, 1'b0, 10'd132},{ 8'd13, 1'b1, 10'd202},
{ 8'd12, 1'b0,  10'd32},{ 8'd12, 1'b0,  10'd72},{ 8'd12, 1'b1, 10'd102},
{ 8'd11, 1'b0,  10'd42},{ 8'd11, 1'b0, 10'd152},{ 8'd11, 1'b1, 10'd192},
{ 8'd10, 1'b0, 10'd122},{ 8'd10, 1'b0, 10'd172},{ 8'd10, 1'b1, 10'd182},
{  8'd9, 1'b0,  10'd43},{  8'd9, 1'b0,  10'd53},{  8'd9, 1'b0, 10'd163},{  8'd9, 1'b1, 10'd173},
{  8'd8, 1'b0,  10'd33},{  8'd8, 1'b0, 10'd143},{  8'd8, 1'b0, 10'd183},{  8'd8, 1'b1, 10'd203},
{  8'd7, 1'b0,  10'd73},{  8'd7, 1'b0,  10'd83},{  8'd7, 1'b0, 10'd123},{  8'd7, 1'b1, 10'd193},
{  8'd6, 1'b0,  10'd13},{  8'd6, 1'b0,  10'd93},{  8'd6, 1'b0, 10'd113},{  8'd6, 1'b1, 10'd133},
{  8'd5, 1'b0,  10'd23},{  8'd5, 1'b0,  10'd63},{  8'd5, 1'b0, 10'd103},{  8'd5, 1'b1, 10'd153},
{  8'd4, 1'b0,  10'd14},{  8'd4, 1'b0,  10'd24},{  8'd4, 1'b0,  10'd34},{  8'd4, 1'b0,  10'd44},{  8'd4, 1'b0,  10'd54},{  8'd4, 1'b0,  10'd64},{  8'd4, 1'b0,  10'd74},{  8'd4, 1'b0,  10'd84},{  8'd4, 1'b0,  10'd94},{  8'd4, 1'b0, 10'd104},{  8'd4, 1'b0, 10'd114},{  8'd4, 1'b0, 10'd124},{  8'd4, 1'b0, 10'd134},{  8'd4, 1'b0, 10'd144},{  8'd4, 1'b0, 10'd154},{  8'd4, 1'b0, 10'd164},{  8'd4, 1'b0, 10'd174},{  8'd4, 1'b0,   10'd4},{  8'd4, 1'b0, 10'd184},{  8'd4, 1'b0, 10'd194},{  8'd4, 1'b1, 10'd204},
{  8'd3, 1'b0,  10'd15},{  8'd3, 1'b0,  10'd25},{  8'd3, 1'b0,  10'd35},{  8'd3, 1'b0,  10'd45},{  8'd3, 1'b0,  10'd55},{  8'd3, 1'b0,  10'd65},{  8'd3, 1'b0,  10'd75},{  8'd3, 1'b0,  10'd85},{  8'd3, 1'b0,  10'd95},{  8'd3, 1'b0, 10'd105},{  8'd3, 1'b0, 10'd115},{  8'd3, 1'b0, 10'd125},{  8'd3, 1'b0, 10'd135},{  8'd3, 1'b0, 10'd145},{  8'd3, 1'b0, 10'd155},{  8'd3, 1'b0, 10'd165},{  8'd3, 1'b0, 10'd175},{  8'd3, 1'b0,   10'd5},{  8'd3, 1'b0, 10'd185},{  8'd3, 1'b0, 10'd195},{  8'd3, 1'b1, 10'd205},
{  8'd2, 1'b0,  10'd16},{  8'd2, 1'b0,  10'd26},{  8'd2, 1'b0,  10'd36},{  8'd2, 1'b0,  10'd46},{  8'd2, 1'b0,  10'd56},{  8'd2, 1'b0,  10'd66},{  8'd2, 1'b0,  10'd76},{  8'd2, 1'b0,  10'd86},{  8'd2, 1'b0,  10'd96},{  8'd2, 1'b0, 10'd106},{  8'd2, 1'b0, 10'd116},{  8'd2, 1'b0, 10'd126},{  8'd2, 1'b0, 10'd136},{  8'd2, 1'b0, 10'd146},{  8'd2, 1'b0, 10'd156},{  8'd2, 1'b0, 10'd166},{  8'd2, 1'b0, 10'd176},{  8'd2, 1'b0,   10'd6},{  8'd2, 1'b0, 10'd186},{  8'd2, 1'b0, 10'd196},{  8'd2, 1'b1, 10'd206},
{  8'd1, 1'b0,  10'd17},{  8'd1, 1'b0,  10'd27},{  8'd1, 1'b0,  10'd37},{  8'd1, 1'b0,  10'd47},{  8'd1, 1'b0,  10'd57},{  8'd1, 1'b0,  10'd67},{  8'd1, 1'b0,  10'd77},{  8'd1, 1'b0,  10'd87},{  8'd1, 1'b0,  10'd97},{  8'd1, 1'b0, 10'd107},{  8'd1, 1'b0, 10'd117},{  8'd1, 1'b0, 10'd127},{  8'd1, 1'b0, 10'd137},{  8'd1, 1'b0, 10'd147},{  8'd1, 1'b0, 10'd157},{  8'd1, 1'b0, 10'd167},{  8'd1, 1'b0, 10'd177},{  8'd1, 1'b0,   10'd7},{  8'd1, 1'b0, 10'd187},{  8'd1, 1'b0, 10'd197},{  8'd1, 1'b1, 10'd207},
{  8'd0, 1'b0,  10'd18},{  8'd0, 1'b0,  10'd28},{  8'd0, 1'b0,  10'd38},{  8'd0, 1'b0,  10'd48},{  8'd0, 1'b0,  10'd58},{  8'd0, 1'b0,  10'd68},{  8'd0, 1'b0,  10'd78},{  8'd0, 1'b0,  10'd88},{  8'd0, 1'b0,  10'd98},{  8'd0, 1'b0, 10'd108},{  8'd0, 1'b0, 10'd118},{  8'd0, 1'b0, 10'd128},{  8'd0, 1'b0, 10'd138},{  8'd0, 1'b0, 10'd148},{  8'd0, 1'b0, 10'd158},{  8'd0, 1'b0, 10'd168},{  8'd0, 1'b0, 10'd178},{  8'd0, 1'b0,   10'd8},{  8'd0, 1'b0, 10'd188},{  8'd0, 1'b0, 10'd198},{  8'd0, 1'b1, 10'd208}
};
localparam int          cSHORT_HS_TAB_26BY45_PACKED_SIZE = 190;
localparam bit [18 : 0] cSHORT_HS_TAB_26BY45_PACKED[cSHORT_HS_TAB_26BY45_PACKED_SIZE] = '{
{  1'b1, 1'b0,  8'd44,    9'd1},{  1'b0, 1'b0,  8'd26,    9'd0},{  1'b0, 1'b0,  8'd13,   9'd39},{  1'b0, 1'b0,   8'd7,  9'd357},{  1'b0, 1'b0,   8'd6,  9'd112},{  1'b0, 1'b0,   8'd5,    9'd0},{  1'b0, 1'b0,   8'd4,   9'd16},{  1'b0, 1'b0,   8'd2,  9'd103},{  1'b0, 1'b0,   8'd1,  9'd323},{  1'b0, 1'b1,   8'd0,   9'd87},
{  1'b0, 1'b0,  8'd27,    9'd0},{  1'b0, 1'b0,  8'd26,    9'd0},{  1'b0, 1'b0,  8'd11,  9'd167},{  1'b0, 1'b0,   8'd7,    9'd0},{  1'b0, 1'b0,   8'd6,  9'd180},{  1'b0, 1'b0,   8'd5,   9'd65},{  1'b0, 1'b0,   8'd4,  9'd347},{  1'b0, 1'b0,   8'd3,   9'd12},{  1'b0, 1'b0,   8'd2,  9'd123},{  1'b0, 1'b1,   8'd0,  9'd114},
{  1'b0, 1'b0,  8'd28,    9'd0},{  1'b0, 1'b0,  8'd27,    9'd0},{  1'b0, 1'b0,  8'd18,  9'd325},{  1'b0, 1'b0,  8'd15,  9'd207},{  1'b0, 1'b0,  8'd11,  9'd269},{  1'b0, 1'b0,   8'd8,  9'd345},{  1'b0, 1'b0,   8'd7,    9'd6},{  1'b0, 1'b0,   8'd4,  9'd151},{  1'b0, 1'b0,   8'd2,  9'd180},{  1'b0, 1'b1,   8'd0,  9'd323},
{  1'b0, 1'b0,  8'd29,    9'd0},{  1'b0, 1'b0,  8'd28,    9'd0},{  1'b0, 1'b0,  8'd22,  9'd219},{  1'b0, 1'b0,  8'd21,    9'd0},{  1'b0, 1'b0,  8'd12,  9'd284},{  1'b0, 1'b0,   8'd9,   9'd44},{  1'b0, 1'b0,   8'd8,  9'd185},{  1'b0, 1'b0,   8'd7,  9'd292},{  1'b0, 1'b0,   8'd6,   9'd80},{  1'b0, 1'b1,   8'd1,  9'd221},
{  1'b0, 1'b0,  8'd30,    9'd0},{  1'b0, 1'b0,  8'd29,    9'd0},{  1'b0, 1'b0,  8'd17,   9'd44},{  1'b0, 1'b0,   8'd7,  9'd177},{  1'b0, 1'b0,   8'd6,  9'd352},{  1'b0, 1'b0,   8'd5,  9'd138},{  1'b0, 1'b0,   8'd4,  9'd266},{  1'b0, 1'b0,   8'd3,   9'd38},{  1'b0, 1'b0,   8'd1,   9'd26},{  1'b0, 1'b1,   8'd0,  9'd355},
{  1'b0, 1'b0,  8'd31,    9'd0},{  1'b0, 1'b0,  8'd30,    9'd0},{  1'b0, 1'b0,  8'd23,   9'd14},{  1'b0, 1'b0,  8'd16,   9'd22},{  1'b0, 1'b0,   8'd7,  9'd118},{  1'b0, 1'b0,   8'd6,  9'd207},{  1'b0, 1'b0,   8'd5,  9'd182},{  1'b0, 1'b0,   8'd3,  9'd140},{  1'b0, 1'b0,   8'd2,  9'd182},{  1'b0, 1'b1,   8'd0,  9'd331},
{  1'b0, 1'b0,  8'd32,    9'd0},{  1'b0, 1'b0,  8'd31,    9'd0},{  1'b0, 1'b0,  8'd19,  9'd215},{  1'b0, 1'b0,  8'd14,   9'd96},{  1'b0, 1'b0,   8'd9,   9'd96},{  1'b0, 1'b0,   8'd7,  9'd263},{  1'b0, 1'b0,   8'd6,   9'd96},{  1'b0, 1'b0,   8'd3,  9'd258},{  1'b0, 1'b0,   8'd2,   9'd11},{  1'b0, 1'b1,   8'd1,  9'd124},
{  1'b0, 1'b0,  8'd33,    9'd0},{  1'b0, 1'b0,  8'd32,    9'd0},{  1'b0, 1'b0,  8'd20,  9'd100},{  1'b0, 1'b0,  8'd12,  9'd131},{  1'b0, 1'b0,   8'd7,  9'd241},{  1'b0, 1'b0,   8'd6,  9'd294},{  1'b0, 1'b0,   8'd5,  9'd116},{  1'b0, 1'b0,   8'd4,  9'd265},{  1'b0, 1'b0,   8'd2,   9'd65},{  1'b0, 1'b1,   8'd0,  9'd321},
{  1'b0, 1'b0,  8'd34,    9'd0},{  1'b0, 1'b0,  8'd33,    9'd0},{  1'b0, 1'b0,  8'd22,   9'd26},{  1'b0, 1'b0,  8'd21,   9'd29},{  1'b0, 1'b0,  8'd20,  9'd318},{  1'b0, 1'b0,  8'd16,  9'd248},{  1'b0, 1'b0,   8'd6,  9'd200},{  1'b0, 1'b0,   8'd4,  9'd303},{  1'b0, 1'b0,   8'd3,  9'd261},{  1'b0, 1'b1,   8'd0,  9'd104},
{  1'b0, 1'b0,  8'd35,    9'd0},{  1'b0, 1'b0,  8'd34,    9'd0},{  1'b0, 1'b0,  8'd25,   9'd50},{  1'b0, 1'b0,  8'd24,  9'd322},{  1'b0, 1'b0,  8'd16,    9'd0},{  1'b0, 1'b0,   8'd6,   9'd72},{  1'b0, 1'b0,   8'd5,  9'd198},{  1'b0, 1'b0,   8'd4,  9'd323},{  1'b0, 1'b0,   8'd2,   9'd72},{  1'b0, 1'b1,   8'd1,   9'd97},
{  1'b0, 1'b0,  8'd36,    9'd0},{  1'b0, 1'b0,  8'd35,    9'd0},{  1'b0, 1'b0,  8'd24,  9'd169},{  1'b0, 1'b0,  8'd23,  9'd292},{  1'b0, 1'b0,  8'd19,  9'd268},{  1'b0, 1'b0,  8'd17,  9'd163},{  1'b0, 1'b0,  8'd13,  9'd149},{  1'b0, 1'b0,   8'd5,  9'd334},{  1'b0, 1'b0,   8'd4,   9'd46},{  1'b0, 1'b1,   8'd1,   9'd66},
{  1'b0, 1'b0,  8'd37,    9'd0},{  1'b0, 1'b0,  8'd36,    9'd0},{  1'b0, 1'b0,  8'd21,   9'd37},{  1'b0, 1'b0,  8'd13,   9'd11},{  1'b0, 1'b0,  8'd12,   9'd68},{  1'b0, 1'b0,   8'd5,  9'd290},{  1'b0, 1'b0,   8'd4,  9'd192},{  1'b0, 1'b0,   8'd3,  9'd304},{  1'b0, 1'b0,   8'd2,  9'd152},{  1'b0, 1'b1,   8'd1,  9'd187},
{  1'b0, 1'b0,  8'd38,    9'd0},{  1'b0, 1'b0,  8'd37,    9'd0},{  1'b0, 1'b0,  8'd23,   9'd53},{  1'b0, 1'b0,  8'd22,  9'd224},{  1'b0, 1'b0,  8'd18,  9'd102},{  1'b0, 1'b0,  8'd10,  9'd313},{  1'b0, 1'b0,   8'd8,  9'd342},{  1'b0, 1'b0,   8'd7,  9'd317},{  1'b0, 1'b0,   8'd1,  9'd145},{  1'b0, 1'b1,   8'd0,  9'd283},
{  1'b0, 1'b0,  8'd39,    9'd0},{  1'b0, 1'b0,  8'd38,    9'd0},{  1'b0, 1'b0,  8'd15,   9'd98},{  1'b0, 1'b0,  8'd14,  9'd220},{  1'b0, 1'b0,   8'd9,  9'd232},{  1'b0, 1'b0,   8'd6,  9'd193},{  1'b0, 1'b0,   8'd4,  9'd136},{  1'b0, 1'b0,   8'd3,  9'd103},{  1'b0, 1'b0,   8'd1,  9'd205},{  1'b0, 1'b1,   8'd0,  9'd201},
{  1'b0, 1'b0,  8'd40,    9'd0},{  1'b0, 1'b0,  8'd39,    9'd0},{  1'b0, 1'b0,  8'd15,   9'd11},{  1'b0, 1'b0,  8'd14,  9'd143},{  1'b0, 1'b0,   8'd7,  9'd192},{  1'b0, 1'b0,   8'd5,  9'd357},{  1'b0, 1'b0,   8'd3,  9'd158},{  1'b0, 1'b0,   8'd2,   9'd13},{  1'b0, 1'b0,   8'd1,   9'd27},{  1'b0, 1'b1,   8'd0,   9'd36},
{  1'b0, 1'b0,  8'd41,    9'd0},{  1'b0, 1'b0,  8'd40,    9'd0},{  1'b0, 1'b0,  8'd10,  9'd323},{  1'b0, 1'b0,   8'd7,  9'd335},{  1'b0, 1'b0,   8'd6,  9'd304},{  1'b0, 1'b0,   8'd5,  9'd221},{  1'b0, 1'b0,   8'd3,  9'd146},{  1'b0, 1'b0,   8'd2,  9'd117},{  1'b0, 1'b0,   8'd1,  9'd173},{  1'b0, 1'b1,   8'd0,  9'd320},
{  1'b0, 1'b0,  8'd42,    9'd0},{  1'b0, 1'b0,  8'd41,    9'd0},{  1'b0, 1'b0,  8'd20,  9'd181},{  1'b0, 1'b0,  8'd18,  9'd339},{  1'b0, 1'b0,  8'd17,  9'd140},{  1'b0, 1'b0,  8'd10,  9'd285},{  1'b0, 1'b0,   8'd5,   9'd44},{  1'b0, 1'b0,   8'd3,  9'd343},{  1'b0, 1'b0,   8'd2,  9'd262},{  1'b0, 1'b1,   8'd0,  9'd321},
{  1'b0, 1'b0,  8'd43,    9'd0},{  1'b0, 1'b0,  8'd42,    9'd0},{  1'b0, 1'b0,  8'd25,  9'd280},{  1'b0, 1'b0,  8'd11,  9'd237},{  1'b0, 1'b0,   8'd6,  9'd182},{  1'b0, 1'b0,   8'd4,   9'd87},{  1'b0, 1'b0,   8'd3,  9'd268},{  1'b0, 1'b0,   8'd2,  9'd103},{  1'b0, 1'b0,   8'd1,  9'd350},{  1'b0, 1'b1,   8'd0,  9'd129},
{  1'b0, 1'b0,  8'd44,    9'd0},{  1'b0, 1'b0,  8'd43,    9'd0},{  1'b0, 1'b0,  8'd25,  9'd143},{  1'b0, 1'b0,  8'd24,   9'd44},{  1'b0, 1'b0,  8'd19,    9'd4},{  1'b0, 1'b0,   8'd7,   9'd39},{  1'b0, 1'b0,   8'd5,  9'd147},{  1'b0, 1'b0,   8'd4,  9'd349},{  1'b0, 1'b0,   8'd3,  9'd278},{  1'b0, 1'b1,   8'd1,  9'd333}
};
localparam bit [18 : 0] cSHORT_HS_V_TAB_26BY45_PACKED[cSHORT_HS_TAB_26BY45_PACKED_SIZE] = '{
{ 8'd44, 1'b0,   10'd0},{ 8'd44, 1'b1, 10'd180},
{ 8'd43, 1'b0, 10'd170},{ 8'd43, 1'b1, 10'd181},
{ 8'd42, 1'b0, 10'd160},{ 8'd42, 1'b1, 10'd171},
{ 8'd41, 1'b0, 10'd150},{ 8'd41, 1'b1, 10'd161},
{ 8'd40, 1'b0, 10'd140},{ 8'd40, 1'b1, 10'd151},
{ 8'd39, 1'b0, 10'd130},{ 8'd39, 1'b1, 10'd141},
{ 8'd38, 1'b0, 10'd120},{ 8'd38, 1'b1, 10'd131},
{ 8'd37, 1'b0, 10'd110},{ 8'd37, 1'b1, 10'd121},
{ 8'd36, 1'b0, 10'd100},{ 8'd36, 1'b1, 10'd111},
{ 8'd35, 1'b0,  10'd90},{ 8'd35, 1'b1, 10'd101},
{ 8'd34, 1'b0,  10'd80},{ 8'd34, 1'b1,  10'd91},
{ 8'd33, 1'b0,  10'd70},{ 8'd33, 1'b1,  10'd81},
{ 8'd32, 1'b0,  10'd60},{ 8'd32, 1'b1,  10'd71},
{ 8'd31, 1'b0,  10'd50},{ 8'd31, 1'b1,  10'd61},
{ 8'd30, 1'b0,  10'd40},{ 8'd30, 1'b1,  10'd51},
{ 8'd29, 1'b0,  10'd30},{ 8'd29, 1'b1,  10'd41},
{ 8'd28, 1'b0,  10'd20},{ 8'd28, 1'b1,  10'd31},
{ 8'd27, 1'b0,  10'd10},{ 8'd27, 1'b1,  10'd21},
{ 8'd26, 1'b0,   10'd1},{ 8'd26, 1'b1,  10'd11},
{ 8'd25, 1'b0,  10'd92},{ 8'd25, 1'b0, 10'd172},{ 8'd25, 1'b1, 10'd182},
{ 8'd24, 1'b0,  10'd93},{ 8'd24, 1'b0, 10'd102},{ 8'd24, 1'b1, 10'd183},
{ 8'd23, 1'b0,  10'd52},{ 8'd23, 1'b0, 10'd103},{ 8'd23, 1'b1, 10'd122},
{ 8'd22, 1'b0,  10'd32},{ 8'd22, 1'b0,  10'd82},{ 8'd22, 1'b1, 10'd123},
{ 8'd21, 1'b0,  10'd33},{ 8'd21, 1'b0,  10'd83},{ 8'd21, 1'b1, 10'd112},
{ 8'd20, 1'b0,  10'd72},{ 8'd20, 1'b0,  10'd84},{ 8'd20, 1'b1, 10'd162},
{ 8'd19, 1'b0,  10'd62},{ 8'd19, 1'b0, 10'd104},{ 8'd19, 1'b1, 10'd184},
{ 8'd18, 1'b0,  10'd22},{ 8'd18, 1'b0, 10'd124},{ 8'd18, 1'b1, 10'd163},
{ 8'd17, 1'b0,  10'd42},{ 8'd17, 1'b0, 10'd105},{ 8'd17, 1'b1, 10'd164},
{ 8'd16, 1'b0,  10'd53},{ 8'd16, 1'b0,  10'd85},{ 8'd16, 1'b1,  10'd94},
{ 8'd15, 1'b0,  10'd23},{ 8'd15, 1'b0, 10'd132},{ 8'd15, 1'b1, 10'd142},
{ 8'd14, 1'b0,  10'd63},{ 8'd14, 1'b0, 10'd133},{ 8'd14, 1'b1, 10'd143},
{ 8'd13, 1'b0,   10'd2},{ 8'd13, 1'b0, 10'd106},{ 8'd13, 1'b1, 10'd113},
{ 8'd12, 1'b0,  10'd34},{ 8'd12, 1'b0,  10'd73},{ 8'd12, 1'b1, 10'd114},
{ 8'd11, 1'b0,  10'd12},{ 8'd11, 1'b0,  10'd24},{ 8'd11, 1'b1, 10'd173},
{ 8'd10, 1'b0, 10'd125},{ 8'd10, 1'b0, 10'd152},{ 8'd10, 1'b1, 10'd165},
{  8'd9, 1'b0,  10'd35},{  8'd9, 1'b0,  10'd64},{  8'd9, 1'b1, 10'd134},
{  8'd8, 1'b0,  10'd25},{  8'd8, 1'b0,  10'd36},{  8'd8, 1'b1, 10'd126},
{  8'd7, 1'b0,   10'd3},{  8'd7, 1'b0,  10'd13},{  8'd7, 1'b0,  10'd26},{  8'd7, 1'b0,  10'd37},{  8'd7, 1'b0,  10'd43},{  8'd7, 1'b0,  10'd54},{  8'd7, 1'b0,  10'd65},{  8'd7, 1'b0,  10'd74},{  8'd7, 1'b0, 10'd127},{  8'd7, 1'b0, 10'd144},{  8'd7, 1'b0, 10'd153},{  8'd7, 1'b1, 10'd185},
{  8'd6, 1'b0,   10'd4},{  8'd6, 1'b0,  10'd14},{  8'd6, 1'b0,  10'd38},{  8'd6, 1'b0,  10'd44},{  8'd6, 1'b0,  10'd55},{  8'd6, 1'b0,  10'd66},{  8'd6, 1'b0,  10'd75},{  8'd6, 1'b0,  10'd86},{  8'd6, 1'b0,  10'd95},{  8'd6, 1'b0, 10'd135},{  8'd6, 1'b0, 10'd154},{  8'd6, 1'b1, 10'd174},
{  8'd5, 1'b0,   10'd5},{  8'd5, 1'b0,  10'd15},{  8'd5, 1'b0,  10'd45},{  8'd5, 1'b0,  10'd56},{  8'd5, 1'b0,  10'd76},{  8'd5, 1'b0,  10'd96},{  8'd5, 1'b0, 10'd107},{  8'd5, 1'b0, 10'd115},{  8'd5, 1'b0, 10'd145},{  8'd5, 1'b0, 10'd155},{  8'd5, 1'b0, 10'd166},{  8'd5, 1'b1, 10'd186},
{  8'd4, 1'b0,   10'd6},{  8'd4, 1'b0,  10'd16},{  8'd4, 1'b0,  10'd27},{  8'd4, 1'b0,  10'd46},{  8'd4, 1'b0,  10'd77},{  8'd4, 1'b0,  10'd87},{  8'd4, 1'b0,  10'd97},{  8'd4, 1'b0, 10'd108},{  8'd4, 1'b0, 10'd116},{  8'd4, 1'b0, 10'd136},{  8'd4, 1'b0, 10'd175},{  8'd4, 1'b1, 10'd187},
{  8'd3, 1'b0,  10'd17},{  8'd3, 1'b0,  10'd47},{  8'd3, 1'b0,  10'd57},{  8'd3, 1'b0,  10'd67},{  8'd3, 1'b0,  10'd88},{  8'd3, 1'b0, 10'd117},{  8'd3, 1'b0, 10'd137},{  8'd3, 1'b0, 10'd146},{  8'd3, 1'b0, 10'd156},{  8'd3, 1'b0, 10'd167},{  8'd3, 1'b0, 10'd176},{  8'd3, 1'b1, 10'd188},
{  8'd2, 1'b0,   10'd7},{  8'd2, 1'b0,  10'd18},{  8'd2, 1'b0,  10'd28},{  8'd2, 1'b0,  10'd58},{  8'd2, 1'b0,  10'd68},{  8'd2, 1'b0,  10'd78},{  8'd2, 1'b0,  10'd98},{  8'd2, 1'b0, 10'd118},{  8'd2, 1'b0, 10'd147},{  8'd2, 1'b0, 10'd157},{  8'd2, 1'b0, 10'd168},{  8'd2, 1'b1, 10'd177},
{  8'd1, 1'b0,   10'd8},{  8'd1, 1'b0,  10'd39},{  8'd1, 1'b0,  10'd48},{  8'd1, 1'b0,  10'd69},{  8'd1, 1'b0,  10'd99},{  8'd1, 1'b0, 10'd109},{  8'd1, 1'b0, 10'd119},{  8'd1, 1'b0, 10'd128},{  8'd1, 1'b0, 10'd138},{  8'd1, 1'b0, 10'd148},{  8'd1, 1'b0, 10'd158},{  8'd1, 1'b0, 10'd178},{  8'd1, 1'b1, 10'd189},
{  8'd0, 1'b0,   10'd9},{  8'd0, 1'b0,  10'd19},{  8'd0, 1'b0,  10'd29},{  8'd0, 1'b0,  10'd49},{  8'd0, 1'b0,  10'd59},{  8'd0, 1'b0,  10'd79},{  8'd0, 1'b0,  10'd89},{  8'd0, 1'b0, 10'd129},{  8'd0, 1'b0, 10'd139},{  8'd0, 1'b0, 10'd149},{  8'd0, 1'b0, 10'd159},{  8'd0, 1'b0, 10'd169},{  8'd0, 1'b1, 10'd179}
};
localparam int          cSHORT_HS_TAB_32BY45_PACKED_SIZE = 169;
localparam bit [18 : 0] cSHORT_HS_TAB_32BY45_PACKED[cSHORT_HS_TAB_32BY45_PACKED_SIZE] = '{
{  1'b1, 1'b0,  8'd44,    9'd1},{  1'b0, 1'b0,  8'd32,    9'd0},{  1'b0, 1'b0,  8'd16,  9'd242},{  1'b0, 1'b0,  8'd15,  9'd254},{  1'b0, 1'b0,  8'd13,   9'd62},{  1'b0, 1'b0,  8'd10,  9'd110},{  1'b0, 1'b0,   8'd9,  9'd149},{  1'b0, 1'b0,   8'd8,  9'd118},{  1'b0, 1'b0,   8'd4,  9'd270},{  1'b0, 1'b0,   8'd3,  9'd199},{  1'b0, 1'b0,   8'd2,   9'd10},{  1'b0, 1'b0,   8'd1,   9'd22},{  1'b0, 1'b1,   8'd0,  9'd324},
{  1'b0, 1'b0,  8'd33,    9'd0},{  1'b0, 1'b0,  8'd32,    9'd0},{  1'b0, 1'b0,  8'd27,  9'd223},{  1'b0, 1'b0,  8'd23,  9'd161},{  1'b0, 1'b0,  8'd21,   9'd43},{  1'b0, 1'b0,  8'd14,  9'd333},{  1'b0, 1'b0,  8'd12,   9'd99},{  1'b0, 1'b0,   8'd6,   9'd83},{  1'b0, 1'b0,   8'd4,  9'd293},{  1'b0, 1'b0,   8'd3,  9'd358},{  1'b0, 1'b0,   8'd2,  9'd223},{  1'b0, 1'b0,   8'd1,  9'd307},{  1'b0, 1'b1,   8'd0,  9'd134},
{  1'b0, 1'b0,  8'd34,    9'd0},{  1'b0, 1'b0,  8'd33,    9'd0},{  1'b0, 1'b0,  8'd31,  9'd117},{  1'b0, 1'b0,  8'd25,  9'd267},{  1'b0, 1'b0,  8'd18,  9'd270},{  1'b0, 1'b0,  8'd17,  9'd139},{  1'b0, 1'b0,  8'd11,  9'd150},{  1'b0, 1'b0,  8'd10,   9'd46},{  1'b0, 1'b0,   8'd4,  9'd189},{  1'b0, 1'b0,   8'd3,  9'd214},{  1'b0, 1'b0,   8'd2,  9'd320},{  1'b0, 1'b0,   8'd1,   9'd24},{  1'b0, 1'b1,   8'd0,   9'd97},
{  1'b0, 1'b0,  8'd35,    9'd0},{  1'b0, 1'b0,  8'd34,    9'd0},{  1'b0, 1'b0,  8'd30,  9'd294},{  1'b0, 1'b0,  8'd23,  9'd137},{  1'b0, 1'b0,  8'd19,   9'd95},{  1'b0, 1'b0,  8'd13,  9'd350},{  1'b0, 1'b0,  8'd12,  9'd240},{  1'b0, 1'b0,   8'd8,  9'd181},{  1'b0, 1'b0,   8'd4,  9'd311},{  1'b0, 1'b0,   8'd3,  9'd325},{  1'b0, 1'b0,   8'd2,  9'd340},{  1'b0, 1'b0,   8'd1,  9'd174},{  1'b0, 1'b1,   8'd0,   9'd14},
{  1'b0, 1'b0,  8'd36,    9'd0},{  1'b0, 1'b0,  8'd35,    9'd0},{  1'b0, 1'b0,  8'd21,  9'd132},{  1'b0, 1'b0,  8'd20,   9'd49},{  1'b0, 1'b0,  8'd19,   9'd19},{  1'b0, 1'b0,  8'd17,   9'd76},{  1'b0, 1'b0,  8'd16,   9'd38},{  1'b0, 1'b0,  8'd15,  9'd351},{  1'b0, 1'b0,  8'd11,  9'd164},{  1'b0, 1'b0,   8'd3,  9'd198},{  1'b0, 1'b0,   8'd2,   9'd64},{  1'b0, 1'b0,   8'd1,  9'd230},{  1'b0, 1'b1,   8'd0,  9'd123},
{  1'b0, 1'b0,  8'd37,    9'd0},{  1'b0, 1'b0,  8'd36,    9'd0},{  1'b0, 1'b0,  8'd28,  9'd156},{  1'b0, 1'b0,  8'd25,  9'd120},{  1'b0, 1'b0,  8'd24,   9'd92},{  1'b0, 1'b0,  8'd22,   9'd69},{  1'b0, 1'b0,   8'd9,  9'd339},{  1'b0, 1'b0,   8'd6,   9'd47},{  1'b0, 1'b0,   8'd4,  9'd350},{  1'b0, 1'b0,   8'd3,   9'd96},{  1'b0, 1'b0,   8'd2,  9'd205},{  1'b0, 1'b0,   8'd1,  9'd195},{  1'b0, 1'b1,   8'd0,   9'd50},
{  1'b0, 1'b0,  8'd38,    9'd0},{  1'b0, 1'b0,  8'd37,    9'd0},{  1'b0, 1'b0,  8'd26,   9'd69},{  1'b0, 1'b0,  8'd24,  9'd240},{  1'b0, 1'b0,  8'd20,  9'd127},{  1'b0, 1'b0,  8'd18,    9'd2},{  1'b0, 1'b0,  8'd12,  9'd231},{  1'b0, 1'b0,   8'd7,  9'd322},{  1'b0, 1'b0,   8'd5,  9'd194},{  1'b0, 1'b0,   8'd4,   9'd26},{  1'b0, 1'b0,   8'd3,  9'd126},{  1'b0, 1'b0,   8'd2,  9'd175},{  1'b0, 1'b1,   8'd0,  9'd273},
{  1'b0, 1'b0,  8'd39,    9'd0},{  1'b0, 1'b0,  8'd38,    9'd0},{  1'b0, 1'b0,  8'd28,  9'd115},{  1'b0, 1'b0,  8'd26,   9'd68},{  1'b0, 1'b0,  8'd23,  9'd307},{  1'b0, 1'b0,  8'd21,  9'd222},{  1'b0, 1'b0,  8'd14,  9'd230},{  1'b0, 1'b0,   8'd9,  9'd209},{  1'b0, 1'b0,   8'd6,   9'd19},{  1'b0, 1'b0,   8'd5,   9'd78},{  1'b0, 1'b0,   8'd4,  9'd327},{  1'b0, 1'b0,   8'd1,  9'd113},{  1'b0, 1'b1,   8'd0,  9'd177},
{  1'b0, 1'b0,  8'd40,    9'd0},{  1'b0, 1'b0,  8'd39,    9'd0},{  1'b0, 1'b0,  8'd29,   9'd95},{  1'b0, 1'b0,  8'd27,  9'd180},{  1'b0, 1'b0,  8'd26,  9'd185},{  1'b0, 1'b0,  8'd19,   9'd34},{  1'b0, 1'b0,  8'd10,  9'd232},{  1'b0, 1'b0,   8'd7,  9'd228},{  1'b0, 1'b0,   8'd4,  9'd335},{  1'b0, 1'b0,   8'd3,  9'd114},{  1'b0, 1'b0,   8'd2,   9'd92},{  1'b0, 1'b0,   8'd1,  9'd212},{  1'b0, 1'b1,   8'd0,  9'd206},
{  1'b0, 1'b0,  8'd41,    9'd0},{  1'b0, 1'b0,  8'd40,    9'd0},{  1'b0, 1'b0,  8'd31,  9'd254},{  1'b0, 1'b0,  8'd30,   9'd23},{  1'b0, 1'b0,  8'd22,  9'd169},{  1'b0, 1'b0,  8'd20,   9'd56},{  1'b0, 1'b0,  8'd15,   9'd53},{  1'b0, 1'b0,   8'd7,  9'd112},{  1'b0, 1'b0,   8'd4,  9'd130},{  1'b0, 1'b0,   8'd3,  9'd343},{  1'b0, 1'b0,   8'd2,  9'd276},{  1'b0, 1'b0,   8'd1,    9'd9},{  1'b0, 1'b1,   8'd0,  9'd213},
{  1'b0, 1'b0,  8'd42,    9'd0},{  1'b0, 1'b0,  8'd41,    9'd0},{  1'b0, 1'b0,  8'd29,   9'd42},{  1'b0, 1'b0,  8'd28,  9'd232},{  1'b0, 1'b0,  8'd25,   9'd58},{  1'b0, 1'b0,  8'd24,  9'd160},{  1'b0, 1'b0,  8'd17,   9'd49},{  1'b0, 1'b0,   8'd5,  9'd166},{  1'b0, 1'b0,   8'd4,  9'd292},{  1'b0, 1'b0,   8'd3,  9'd280},{  1'b0, 1'b0,   8'd2,  9'd215},{  1'b0, 1'b0,   8'd1,  9'd350},{  1'b0, 1'b1,   8'd0,   9'd47},
{  1'b0, 1'b0,  8'd43,    9'd0},{  1'b0, 1'b0,  8'd42,    9'd0},{  1'b0, 1'b0,  8'd27,  9'd175},{  1'b0, 1'b0,  8'd18,  9'd330},{  1'b0, 1'b0,  8'd16,  9'd181},{  1'b0, 1'b0,  8'd13,  9'd176},{  1'b0, 1'b0,  8'd11,  9'd274},{  1'b0, 1'b0,   8'd5,  9'd210},{  1'b0, 1'b0,   8'd4,  9'd312},{  1'b0, 1'b0,   8'd3,  9'd234},{  1'b0, 1'b0,   8'd2,  9'd276},{  1'b0, 1'b0,   8'd1,  9'd218},{  1'b0, 1'b1,   8'd0,   9'd25},
{  1'b0, 1'b0,  8'd44,    9'd0},{  1'b0, 1'b0,  8'd43,    9'd0},{  1'b0, 1'b0,  8'd31,   9'd29},{  1'b0, 1'b0,  8'd30,  9'd170},{  1'b0, 1'b0,  8'd29,  9'd184},{  1'b0, 1'b0,  8'd22,  9'd129},{  1'b0, 1'b0,  8'd14,   9'd30},{  1'b0, 1'b0,   8'd8,  9'd228},{  1'b0, 1'b0,   8'd5,  9'd216},{  1'b0, 1'b0,   8'd4,  9'd255},{  1'b0, 1'b0,   8'd3,  9'd144},{  1'b0, 1'b0,   8'd2,  9'd212},{  1'b0, 1'b1,   8'd1,  9'd199}
};
localparam bit [18 : 0] cSHORT_HS_V_TAB_32BY45_PACKED[cSHORT_HS_TAB_32BY45_PACKED_SIZE] = '{
{ 8'd44, 1'b0,   10'd0},{ 8'd44, 1'b1, 10'd156},
{ 8'd43, 1'b0, 10'd143},{ 8'd43, 1'b1, 10'd157},
{ 8'd42, 1'b0, 10'd130},{ 8'd42, 1'b1, 10'd144},
{ 8'd41, 1'b0, 10'd117},{ 8'd41, 1'b1, 10'd131},
{ 8'd40, 1'b0, 10'd104},{ 8'd40, 1'b1, 10'd118},
{ 8'd39, 1'b0,  10'd91},{ 8'd39, 1'b1, 10'd105},
{ 8'd38, 1'b0,  10'd78},{ 8'd38, 1'b1,  10'd92},
{ 8'd37, 1'b0,  10'd65},{ 8'd37, 1'b1,  10'd79},
{ 8'd36, 1'b0,  10'd52},{ 8'd36, 1'b1,  10'd66},
{ 8'd35, 1'b0,  10'd39},{ 8'd35, 1'b1,  10'd53},
{ 8'd34, 1'b0,  10'd26},{ 8'd34, 1'b1,  10'd40},
{ 8'd33, 1'b0,  10'd13},{ 8'd33, 1'b1,  10'd27},
{ 8'd32, 1'b0,   10'd1},{ 8'd32, 1'b1,  10'd14},
{ 8'd31, 1'b0,  10'd28},{ 8'd31, 1'b0, 10'd119},{ 8'd31, 1'b1, 10'd158},
{ 8'd30, 1'b0,  10'd41},{ 8'd30, 1'b0, 10'd120},{ 8'd30, 1'b1, 10'd159},
{ 8'd29, 1'b0, 10'd106},{ 8'd29, 1'b0, 10'd132},{ 8'd29, 1'b1, 10'd160},
{ 8'd28, 1'b0,  10'd67},{ 8'd28, 1'b0,  10'd93},{ 8'd28, 1'b1, 10'd133},
{ 8'd27, 1'b0,  10'd15},{ 8'd27, 1'b0, 10'd107},{ 8'd27, 1'b1, 10'd145},
{ 8'd26, 1'b0,  10'd80},{ 8'd26, 1'b0,  10'd94},{ 8'd26, 1'b1, 10'd108},
{ 8'd25, 1'b0,  10'd29},{ 8'd25, 1'b0,  10'd68},{ 8'd25, 1'b1, 10'd134},
{ 8'd24, 1'b0,  10'd69},{ 8'd24, 1'b0,  10'd81},{ 8'd24, 1'b1, 10'd135},
{ 8'd23, 1'b0,  10'd16},{ 8'd23, 1'b0,  10'd42},{ 8'd23, 1'b1,  10'd95},
{ 8'd22, 1'b0,  10'd70},{ 8'd22, 1'b0, 10'd121},{ 8'd22, 1'b1, 10'd161},
{ 8'd21, 1'b0,  10'd17},{ 8'd21, 1'b0,  10'd54},{ 8'd21, 1'b1,  10'd96},
{ 8'd20, 1'b0,  10'd55},{ 8'd20, 1'b0,  10'd82},{ 8'd20, 1'b1, 10'd122},
{ 8'd19, 1'b0,  10'd43},{ 8'd19, 1'b0,  10'd56},{ 8'd19, 1'b1, 10'd109},
{ 8'd18, 1'b0,  10'd30},{ 8'd18, 1'b0,  10'd83},{ 8'd18, 1'b1, 10'd146},
{ 8'd17, 1'b0,  10'd31},{ 8'd17, 1'b0,  10'd57},{ 8'd17, 1'b1, 10'd136},
{ 8'd16, 1'b0,   10'd2},{ 8'd16, 1'b0,  10'd58},{ 8'd16, 1'b1, 10'd147},
{ 8'd15, 1'b0,   10'd3},{ 8'd15, 1'b0,  10'd59},{ 8'd15, 1'b1, 10'd123},
{ 8'd14, 1'b0,  10'd18},{ 8'd14, 1'b0,  10'd97},{ 8'd14, 1'b1, 10'd162},
{ 8'd13, 1'b0,   10'd4},{ 8'd13, 1'b0,  10'd44},{ 8'd13, 1'b1, 10'd148},
{ 8'd12, 1'b0,  10'd19},{ 8'd12, 1'b0,  10'd45},{ 8'd12, 1'b1,  10'd84},
{ 8'd11, 1'b0,  10'd32},{ 8'd11, 1'b0,  10'd60},{ 8'd11, 1'b1, 10'd149},
{ 8'd10, 1'b0,   10'd5},{ 8'd10, 1'b0,  10'd33},{ 8'd10, 1'b1, 10'd110},
{  8'd9, 1'b0,   10'd6},{  8'd9, 1'b0,  10'd71},{  8'd9, 1'b1,  10'd98},
{  8'd8, 1'b0,   10'd7},{  8'd8, 1'b0,  10'd46},{  8'd8, 1'b1, 10'd163},
{  8'd7, 1'b0,  10'd85},{  8'd7, 1'b0, 10'd111},{  8'd7, 1'b1, 10'd124},
{  8'd6, 1'b0,  10'd20},{  8'd6, 1'b0,  10'd72},{  8'd6, 1'b1,  10'd99},
{  8'd5, 1'b0,  10'd86},{  8'd5, 1'b0, 10'd100},{  8'd5, 1'b0, 10'd137},{  8'd5, 1'b0, 10'd150},{  8'd5, 1'b1, 10'd164},
{  8'd4, 1'b0,   10'd8},{  8'd4, 1'b0,  10'd21},{  8'd4, 1'b0,  10'd34},{  8'd4, 1'b0,  10'd47},{  8'd4, 1'b0,  10'd73},{  8'd4, 1'b0,  10'd87},{  8'd4, 1'b0, 10'd101},{  8'd4, 1'b0, 10'd112},{  8'd4, 1'b0, 10'd125},{  8'd4, 1'b0, 10'd138},{  8'd4, 1'b0, 10'd151},{  8'd4, 1'b1, 10'd165},
{  8'd3, 1'b0,   10'd9},{  8'd3, 1'b0,  10'd22},{  8'd3, 1'b0,  10'd35},{  8'd3, 1'b0,  10'd48},{  8'd3, 1'b0,  10'd61},{  8'd3, 1'b0,  10'd74},{  8'd3, 1'b0,  10'd88},{  8'd3, 1'b0, 10'd113},{  8'd3, 1'b0, 10'd126},{  8'd3, 1'b0, 10'd139},{  8'd3, 1'b0, 10'd152},{  8'd3, 1'b1, 10'd166},
{  8'd2, 1'b0,  10'd10},{  8'd2, 1'b0,  10'd23},{  8'd2, 1'b0,  10'd36},{  8'd2, 1'b0,  10'd49},{  8'd2, 1'b0,  10'd62},{  8'd2, 1'b0,  10'd75},{  8'd2, 1'b0,  10'd89},{  8'd2, 1'b0, 10'd114},{  8'd2, 1'b0, 10'd127},{  8'd2, 1'b0, 10'd140},{  8'd2, 1'b0, 10'd153},{  8'd2, 1'b1, 10'd167},
{  8'd1, 1'b0,  10'd11},{  8'd1, 1'b0,  10'd24},{  8'd1, 1'b0,  10'd37},{  8'd1, 1'b0,  10'd50},{  8'd1, 1'b0,  10'd63},{  8'd1, 1'b0,  10'd76},{  8'd1, 1'b0, 10'd102},{  8'd1, 1'b0, 10'd115},{  8'd1, 1'b0, 10'd128},{  8'd1, 1'b0, 10'd141},{  8'd1, 1'b0, 10'd154},{  8'd1, 1'b1, 10'd168},
{  8'd0, 1'b0,  10'd12},{  8'd0, 1'b0,  10'd25},{  8'd0, 1'b0,  10'd38},{  8'd0, 1'b0,  10'd51},{  8'd0, 1'b0,  10'd64},{  8'd0, 1'b0,  10'd77},{  8'd0, 1'b0,  10'd90},{  8'd0, 1'b0, 10'd103},{  8'd0, 1'b0, 10'd116},{  8'd0, 1'b0, 10'd129},{  8'd0, 1'b0, 10'd142},{  8'd0, 1'b1, 10'd155}
};
