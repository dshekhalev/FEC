//
// (!!!) IT'S GENERATED short table for cCODE_5by6 coderate, 2304 bits do 8 LLR per cycle(!!!)
//
  addr_tab[0][0][0] = '{baddr:1, offset:'{0, 511, 511, 511, 511, 511, 511, 511}, offsetm:'{0, 511, 511, 511, 511, 511, 511, 511}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}, invsela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[0][1][0] = '{baddr:4, offset:'{0, 511, 511, 511, 511, 511, 511, 511}, offsetm:'{0, 511, 511, 511, 511, 511, 511, 511}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}, invsela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[0][2][0] = '{baddr:7, offset:'{0, 0, 0, 0, 0, 0, 0, 511}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 511}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}, invsela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[0][3][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[0][4][0] = '{baddr:6, offset:'{0, 0, 0, 0, 0, 0, 0, 511}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 511}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}, invsela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[0][5][0] = '{baddr:1, offset:'{0, 0, 0, 0, 511, 511, 511, 511}, offsetm:'{0, 0, 0, 0, 511, 511, 511, 511}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}, invsela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[0][6][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[0][7][0] = '{baddr:0, offset:'{0, 0, 0, 11, 11, 11, 11, 11}, offsetm:'{0, 0, 0, 511, 511, 511, 511, 511}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}, invsela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[0][8][0] = '{baddr:11, offset:'{0, 0, 0, 0, 511, 511, 511, 511}, offsetm:'{0, 0, 0, 0, 511, 511, 511, 511}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}, invsela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[0][9][0] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[0][10][0] = '{baddr:11, offset:'{0, 0, 0, 0, 0, 0, 511, 511}, offsetm:'{0, 0, 0, 0, 0, 0, 511, 511}, sela:'{6, 7, 0, 1, 2, 3, 4, 5}, invsela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[0][11][0] = '{baddr:7, offset:'{0, 0, 0, 0, 511, 511, 511, 511}, offsetm:'{0, 0, 0, 0, 511, 511, 511, 511}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}, invsela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[0][12][0] = '{baddr:11, offset:'{0, 0, 511, 511, 511, 511, 511, 511}, offsetm:'{0, 0, 511, 511, 511, 511, 511, 511}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}, invsela:'{6, 7, 0, 1, 2, 3, 4, 5}};
  addr_tab[0][13][0] = '{baddr:5, offset:'{0, 511, 511, 511, 511, 511, 511, 511}, offsetm:'{0, 511, 511, 511, 511, 511, 511, 511}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}, invsela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[0][14][0] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 511, 511, 511}, offsetm:'{0, 0, 0, 0, 0, 511, 511, 511}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}, invsela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[0][15][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[0][16][0] = '{baddr:5, offset:'{0, 0, 0, 0, 511, 511, 511, 511}, offsetm:'{0, 0, 0, 0, 511, 511, 511, 511}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}, invsela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[0][17][0] = '{baddr:3, offset:'{0, 0, 0, 0, 511, 511, 511, 511}, offsetm:'{0, 0, 0, 0, 511, 511, 511, 511}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}, invsela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[0][18][0] = '{baddr:1, offset:'{0, 0, 0, 0, 511, 511, 511, 511}, offsetm:'{0, 0, 0, 0, 511, 511, 511, 511}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}, invsela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[0][19][0] = '{baddr:10, offset:'{0, 0, 0, 0, 0, 511, 511, 511}, offsetm:'{0, 0, 0, 0, 0, 511, 511, 511}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}, invsela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[0][20][0] = '{baddr:10, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[0][21][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[0][22][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[0][23][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[1][0][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[1][1][0] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 511, 511}, offsetm:'{0, 0, 0, 0, 0, 0, 511, 511}, sela:'{6, 7, 0, 1, 2, 3, 4, 5}, invsela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[1][2][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[1][3][0] = '{baddr:5, offset:'{0, 0, 0, 0, 511, 511, 511, 511}, offsetm:'{0, 0, 0, 0, 511, 511, 511, 511}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}, invsela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[1][4][0] = '{baddr:5, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[1][5][0] = '{baddr:6, offset:'{0, 0, 0, 0, 0, 0, 0, 511}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 511}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}, invsela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[1][6][0] = '{baddr:2, offset:'{0, 0, 0, 0, 511, 511, 511, 511}, offsetm:'{0, 0, 0, 0, 511, 511, 511, 511}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}, invsela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[1][7][0] = '{baddr:10, offset:'{0, 0, 0, 0, 0, 0, 0, 511}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 511}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}, invsela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[1][8][0] = '{baddr:6, offset:'{0, 0, 0, 0, 0, 0, 0, 511}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 511}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}, invsela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[1][9][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[1][10][0] = '{baddr:6, offset:'{0, 511, 511, 511, 511, 511, 511, 511}, offsetm:'{0, 511, 511, 511, 511, 511, 511, 511}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}, invsela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[1][11][0] = '{baddr:3, offset:'{0, 0, 0, 0, 0, 511, 511, 511}, offsetm:'{0, 0, 0, 0, 0, 511, 511, 511}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}, invsela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[1][12][0] = '{baddr:2, offset:'{0, 0, 0, 0, 511, 511, 511, 511}, offsetm:'{0, 0, 0, 0, 511, 511, 511, 511}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}, invsela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[1][13][0] = '{baddr:9, offset:'{0, 0, 0, 0, 0, 0, 0, 511}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 511}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}, invsela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[1][14][0] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 511, 511}, offsetm:'{0, 0, 0, 0, 0, 0, 511, 511}, sela:'{6, 7, 0, 1, 2, 3, 4, 5}, invsela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[1][15][0] = '{baddr:9, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[1][16][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[1][17][0] = '{baddr:6, offset:'{0, 0, 0, 0, 511, 511, 511, 511}, offsetm:'{0, 0, 0, 0, 511, 511, 511, 511}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}, invsela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[1][18][0] = '{baddr:7, offset:'{0, 511, 511, 511, 511, 511, 511, 511}, offsetm:'{0, 511, 511, 511, 511, 511, 511, 511}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}, invsela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[1][19][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[1][20][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[1][21][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[1][22][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[1][23][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[2][0][0] = '{baddr:7, offset:'{0, 0, 0, 511, 511, 511, 511, 511}, offsetm:'{0, 0, 0, 511, 511, 511, 511, 511}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}, invsela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[2][1][0] = '{baddr:11, offset:'{0, 511, 511, 511, 511, 511, 511, 511}, offsetm:'{0, 511, 511, 511, 511, 511, 511, 511}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}, invsela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[2][2][0] = '{baddr:11, offset:'{0, 0, 0, 511, 511, 511, 511, 511}, offsetm:'{0, 0, 0, 511, 511, 511, 511, 511}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}, invsela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[2][3][0] = '{baddr:1, offset:'{0, 0, 0, 0, 511, 511, 511, 511}, offsetm:'{0, 0, 0, 0, 511, 511, 511, 511}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}, invsela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[2][4][0] = '{baddr:9, offset:'{0, 0, 0, 511, 511, 511, 511, 511}, offsetm:'{0, 0, 0, 511, 511, 511, 511, 511}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}, invsela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[2][5][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[2][6][0] = '{baddr:3, offset:'{0, 0, 0, 0, 0, 511, 511, 511}, offsetm:'{0, 0, 0, 0, 0, 511, 511, 511}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}, invsela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[2][7][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[2][8][0] = '{baddr:4, offset:'{0, 0, 0, 0, 0, 0, 0, 511}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 511}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}, invsela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[2][9][0] = '{baddr:3, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[2][10][0] = '{baddr:0, offset:'{0, 0, 0, 11, 11, 11, 11, 11}, offsetm:'{0, 0, 0, 511, 511, 511, 511, 511}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}, invsela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[2][11][0] = '{baddr:8, offset:'{0, 0, 0, 0, 0, 511, 511, 511}, offsetm:'{0, 0, 0, 0, 0, 511, 511, 511}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}, invsela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[2][12][0] = '{baddr:11, offset:'{0, 511, 511, 511, 511, 511, 511, 511}, offsetm:'{0, 511, 511, 511, 511, 511, 511, 511}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}, invsela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[2][13][0] = '{baddr:2, offset:'{0, 511, 511, 511, 511, 511, 511, 511}, offsetm:'{0, 511, 511, 511, 511, 511, 511, 511}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}, invsela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[2][14][0] = '{baddr:11, offset:'{0, 0, 0, 0, 0, 0, 511, 511}, offsetm:'{0, 0, 0, 0, 0, 0, 511, 511}, sela:'{6, 7, 0, 1, 2, 3, 4, 5}, invsela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[2][15][0] = '{baddr:10, offset:'{0, 0, 0, 0, 0, 0, 511, 511}, offsetm:'{0, 0, 0, 0, 0, 0, 511, 511}, sela:'{6, 7, 0, 1, 2, 3, 4, 5}, invsela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[2][16][0] = '{baddr:8, offset:'{0, 0, 0, 0, 511, 511, 511, 511}, offsetm:'{0, 0, 0, 0, 511, 511, 511, 511}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}, invsela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[2][17][0] = '{baddr:11, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[2][18][0] = '{baddr:9, offset:'{0, 0, 0, 511, 511, 511, 511, 511}, offsetm:'{0, 0, 0, 511, 511, 511, 511, 511}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}, invsela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[2][19][0] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 511}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 511}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}, invsela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[2][20][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[2][21][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[2][22][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[2][23][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[3][0][0] = '{baddr:9, offset:'{0, 0, 0, 0, 511, 511, 511, 511}, offsetm:'{0, 0, 0, 0, 511, 511, 511, 511}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}, invsela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[3][1][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[3][2][0] = '{baddr:7, offset:'{0, 0, 511, 511, 511, 511, 511, 511}, offsetm:'{0, 0, 511, 511, 511, 511, 511, 511}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}, invsela:'{6, 7, 0, 1, 2, 3, 4, 5}};
  addr_tab[3][3][0] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 511}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 511}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}, invsela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[3][4][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[3][5][0] = '{baddr:5, offset:'{0, 0, 0, 0, 511, 511, 511, 511}, offsetm:'{0, 0, 0, 0, 511, 511, 511, 511}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}, invsela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[3][6][0] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 511, 511, 511}, offsetm:'{0, 0, 0, 0, 0, 511, 511, 511}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}, invsela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[3][7][0] = '{baddr:2, offset:'{0, 0, 511, 511, 511, 511, 511, 511}, offsetm:'{0, 0, 511, 511, 511, 511, 511, 511}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}, invsela:'{6, 7, 0, 1, 2, 3, 4, 5}};
  addr_tab[3][8][0] = '{baddr:2, offset:'{0, 0, 0, 511, 511, 511, 511, 511}, offsetm:'{0, 0, 0, 511, 511, 511, 511, 511}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}, invsela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[3][9][0] = '{baddr:3, offset:'{0, 0, 0, 0, 511, 511, 511, 511}, offsetm:'{0, 0, 0, 0, 511, 511, 511, 511}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}, invsela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[3][10][0] = '{baddr:7, offset:'{0, 0, 0, 0, 0, 511, 511, 511}, offsetm:'{0, 0, 0, 0, 0, 511, 511, 511}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}, invsela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[3][11][0] = '{baddr:0, offset:'{0, 0, 11, 11, 11, 11, 11, 11}, offsetm:'{0, 0, 511, 511, 511, 511, 511, 511}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}, invsela:'{6, 7, 0, 1, 2, 3, 4, 5}};
  addr_tab[3][12][0] = '{baddr:4, offset:'{0, 0, 0, 0, 0, 511, 511, 511}, offsetm:'{0, 0, 0, 0, 0, 511, 511, 511}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}, invsela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[3][13][0] = '{baddr:0, offset:'{0, 0, 0, 0, 11, 11, 11, 11}, offsetm:'{0, 0, 0, 0, 511, 511, 511, 511}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}, invsela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[3][14][0] = '{baddr:8, offset:'{0, 511, 511, 511, 511, 511, 511, 511}, offsetm:'{0, 511, 511, 511, 511, 511, 511, 511}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}, invsela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[3][15][0] = '{baddr:4, offset:'{0, 0, 0, 0, 0, 0, 511, 511}, offsetm:'{0, 0, 0, 0, 0, 0, 511, 511}, sela:'{6, 7, 0, 1, 2, 3, 4, 5}, invsela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[3][16][0] = '{baddr:11, offset:'{0, 0, 0, 0, 511, 511, 511, 511}, offsetm:'{0, 0, 0, 0, 511, 511, 511, 511}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}, invsela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[3][17][0] = '{baddr:0, offset:'{0, 0, 0, 0, 11, 11, 11, 11}, offsetm:'{0, 0, 0, 0, 511, 511, 511, 511}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}, invsela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[3][18][0] = '{baddr:2, offset:'{0, 0, 0, 511, 511, 511, 511, 511}, offsetm:'{0, 0, 0, 511, 511, 511, 511, 511}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}, invsela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[3][19][0] = '{baddr:9, offset:'{0, 0, 511, 511, 511, 511, 511, 511}, offsetm:'{0, 0, 511, 511, 511, 511, 511, 511}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}, invsela:'{6, 7, 0, 1, 2, 3, 4, 5}};
  addr_tab[3][20][0] = '{baddr:10, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[3][21][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[3][22][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[3][23][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}, invsela:'{0, 1, 2, 3, 4, 5, 6, 7}};
