localparam int          cLARGE_HS_TAB_1BY4_PACKED_SIZE = 540;
localparam bit [18 : 0] cLARGE_HS_TAB_1BY4_PACKED[cLARGE_HS_TAB_1BY4_PACKED_SIZE] = '{
{  1'b1, 1'b0, 8'd179,    9'd1},{  1'b0, 1'b0,  8'd45,    9'd0},{  1'b0, 1'b0,  8'd27,   9'd69},{  1'b0, 1'b1,   8'd0,    9'd4},
{  1'b0, 1'b0,  8'd46,    9'd0},{  1'b0, 1'b0,  8'd45,    9'd0},{  1'b0, 1'b0,  8'd44,  9'd243},{  1'b0, 1'b1,  8'd28,  9'd267},
{  1'b0, 1'b0,  8'd47,    9'd0},{  1'b0, 1'b0,  8'd46,    9'd0},{  1'b0, 1'b0,  8'd14,   9'd20},{  1'b0, 1'b1,   8'd6,   9'd14},
{  1'b0, 1'b0,  8'd48,    9'd0},{  1'b0, 1'b0,  8'd47,    9'd0},{  1'b0, 1'b0,  8'd20,  9'd325},{  1'b0, 1'b1,  8'd13,  9'd332},
{  1'b0, 1'b0,  8'd49,    9'd0},{  1'b0, 1'b0,  8'd48,    9'd0},{  1'b0, 1'b0,  8'd11,  9'd355},{  1'b0, 1'b1,   8'd1,  9'd123},
{  1'b0, 1'b0,  8'd50,    9'd0},{  1'b0, 1'b0,  8'd49,    9'd0},{  1'b0, 1'b0,  8'd25,  9'd325},{  1'b0, 1'b1,   8'd4,  9'd201},
{  1'b0, 1'b0,  8'd51,    9'd0},{  1'b0, 1'b0,  8'd50,    9'd0},{  1'b0, 1'b0,   8'd5,  9'd103},{  1'b0, 1'b1,   8'd5,  9'd189},
{  1'b0, 1'b0,  8'd52,    9'd0},{  1'b0, 1'b0,  8'd51,    9'd0},{  1'b0, 1'b0,  8'd12,  9'd311},{  1'b0, 1'b1,  8'd10,  9'd101},
{  1'b0, 1'b0,  8'd53,    9'd0},{  1'b0, 1'b0,  8'd52,    9'd0},{  1'b0, 1'b0,  8'd35,  9'd226},{  1'b0, 1'b1,  8'd24,  9'd286},
{  1'b0, 1'b0,  8'd54,    9'd0},{  1'b0, 1'b0,  8'd53,    9'd0},{  1'b0, 1'b0,  8'd41,  9'd219},{  1'b0, 1'b1,  8'd17,   9'd47},
{  1'b0, 1'b0,  8'd55,    9'd0},{  1'b0, 1'b0,  8'd54,    9'd0},{  1'b0, 1'b0,  8'd10,   9'd63},{  1'b0, 1'b1,   8'd9,  9'd312},
{  1'b0, 1'b0,  8'd56,    9'd0},{  1'b0, 1'b0,  8'd55,    9'd0},{  1'b0, 1'b0,  8'd12,   9'd62},{  1'b0, 1'b1,   8'd2,   9'd97},
{  1'b0, 1'b0,  8'd57,    9'd0},{  1'b0, 1'b0,  8'd56,    9'd0},{  1'b0, 1'b0,  8'd15,  9'd164},{  1'b0, 1'b1,   8'd8,  9'd223},
{  1'b0, 1'b0,  8'd58,    9'd0},{  1'b0, 1'b0,  8'd57,    9'd0},{  1'b0, 1'b0,  8'd42,  9'd243},{  1'b0, 1'b1,  8'd14,  9'd237},
{  1'b0, 1'b0,  8'd59,    9'd0},{  1'b0, 1'b0,  8'd58,    9'd0},{  1'b0, 1'b0,  8'd29,   9'd54},{  1'b0, 1'b1,  8'd11,  9'd144},
{  1'b0, 1'b0,  8'd60,    9'd0},{  1'b0, 1'b0,  8'd59,    9'd0},{  1'b0, 1'b0,   8'd2,  9'd224},{  1'b0, 1'b1,   8'd0,  9'd137},
{  1'b0, 1'b0,  8'd61,    9'd0},{  1'b0, 1'b0,  8'd60,    9'd0},{  1'b0, 1'b0,   8'd7,  9'd328},{  1'b0, 1'b1,   8'd0,   9'd46},
{  1'b0, 1'b0,  8'd62,    9'd0},{  1'b0, 1'b0,  8'd61,    9'd0},{  1'b0, 1'b0,  8'd12,   9'd92},{  1'b0, 1'b1,   8'd8,  9'd324},
{  1'b0, 1'b0,  8'd63,    9'd0},{  1'b0, 1'b0,  8'd62,    9'd0},{  1'b0, 1'b0,  8'd40,  9'd126},{  1'b0, 1'b1,   8'd9,  9'd206},
{  1'b0, 1'b0,  8'd64,    9'd0},{  1'b0, 1'b0,  8'd63,    9'd0},{  1'b0, 1'b0,  8'd12,  9'd195},{  1'b0, 1'b1,   8'd8,  9'd309},
{  1'b0, 1'b0,  8'd65,    9'd0},{  1'b0, 1'b0,  8'd64,    9'd0},{  1'b0, 1'b0,  8'd30,   9'd96},{  1'b0, 1'b1,  8'd11,  9'd326},
{  1'b0, 1'b0,  8'd66,    9'd0},{  1'b0, 1'b0,  8'd65,    9'd0},{  1'b0, 1'b0,  8'd23,  9'd179},{  1'b0, 1'b1,  8'd14,  9'd203},
{  1'b0, 1'b0,  8'd67,    9'd0},{  1'b0, 1'b0,  8'd66,    9'd0},{  1'b0, 1'b0,  8'd35,  9'd273},{  1'b0, 1'b1,   8'd1,  9'd185},
{  1'b0, 1'b0,  8'd68,    9'd0},{  1'b0, 1'b0,  8'd67,    9'd0},{  1'b0, 1'b0,  8'd36,   9'd56},{  1'b0, 1'b1,  8'd10,  9'd192},
{  1'b0, 1'b0,  8'd69,    9'd0},{  1'b0, 1'b0,  8'd68,    9'd0},{  1'b0, 1'b0,   8'd8,  9'd214},{  1'b0, 1'b1,   8'd6,  9'd333},
{  1'b0, 1'b0,  8'd70,    9'd0},{  1'b0, 1'b0,  8'd69,    9'd0},{  1'b0, 1'b0,  8'd13,  9'd277},{  1'b0, 1'b1,   8'd5,  9'd166},
{  1'b0, 1'b0,  8'd71,    9'd0},{  1'b0, 1'b0,  8'd70,    9'd0},{  1'b0, 1'b0,  8'd34,  9'd181},{  1'b0, 1'b1,  8'd17,  9'd259},
{  1'b0, 1'b0,  8'd72,    9'd0},{  1'b0, 1'b0,  8'd71,    9'd0},{  1'b0, 1'b0,   8'd4,  9'd213},{  1'b0, 1'b1,   8'd3,   9'd66},
{  1'b0, 1'b0,  8'd73,    9'd0},{  1'b0, 1'b0,  8'd72,    9'd0},{  1'b0, 1'b0,  8'd14,  9'd287},{  1'b0, 1'b1,   8'd7,  9'd298},
{  1'b0, 1'b0,  8'd74,    9'd0},{  1'b0, 1'b0,  8'd73,    9'd0},{  1'b0, 1'b0,   8'd2,  9'd107},{  1'b0, 1'b1,   8'd0,  9'd311},
{  1'b0, 1'b0,  8'd75,    9'd0},{  1'b0, 1'b0,  8'd74,    9'd0},{  1'b0, 1'b0,  8'd30,  9'd125},{  1'b0, 1'b1,   8'd6,  9'd312},
{  1'b0, 1'b0,  8'd76,    9'd0},{  1'b0, 1'b0,  8'd75,    9'd0},{  1'b0, 1'b0,   8'd5,  9'd242},{  1'b0, 1'b1,   8'd4,   9'd74},
{  1'b0, 1'b0,  8'd77,    9'd0},{  1'b0, 1'b0,  8'd76,    9'd0},{  1'b0, 1'b0,  8'd36,  9'd180},{  1'b0, 1'b1,  8'd24,  9'd229},
{  1'b0, 1'b0,  8'd78,    9'd0},{  1'b0, 1'b0,  8'd77,    9'd0},{  1'b0, 1'b0,  8'd25,  9'd263},{  1'b0, 1'b1,  8'd11,  9'd180},
{  1'b0, 1'b0,  8'd79,    9'd0},{  1'b0, 1'b0,  8'd78,    9'd0},{  1'b0, 1'b0,   8'd8,  9'd160},{  1'b0, 1'b1,   8'd1,  9'd274},
{  1'b0, 1'b0,  8'd80,    9'd0},{  1'b0, 1'b0,  8'd79,    9'd0},{  1'b0, 1'b0,  8'd40,   9'd69},{  1'b0, 1'b1,  8'd10,  9'd229},
{  1'b0, 1'b0,  8'd81,    9'd0},{  1'b0, 1'b0,  8'd80,    9'd0},{  1'b0, 1'b0,   8'd6,  9'd171},{  1'b0, 1'b1,   8'd4,  9'd299},
{  1'b0, 1'b0,  8'd82,    9'd0},{  1'b0, 1'b0,  8'd81,    9'd0},{  1'b0, 1'b0,   8'd9,  9'd253},{  1'b0, 1'b1,   8'd1,  9'd153},
{  1'b0, 1'b0,  8'd83,    9'd0},{  1'b0, 1'b0,  8'd82,    9'd0},{  1'b0, 1'b0,  8'd27,  9'd162},{  1'b0, 1'b1,   8'd3,  9'd296},
{  1'b0, 1'b0,  8'd84,    9'd0},{  1'b0, 1'b0,  8'd83,    9'd0},{  1'b0, 1'b0,  8'd19,  9'd106},{  1'b0, 1'b1,   8'd9,   9'd33},
{  1'b0, 1'b0,  8'd85,    9'd0},{  1'b0, 1'b0,  8'd84,    9'd0},{  1'b0, 1'b0,  8'd33,   9'd65},{  1'b0, 1'b1,   8'd5,  9'd300},
{  1'b0, 1'b0,  8'd86,    9'd0},{  1'b0, 1'b0,  8'd85,    9'd0},{  1'b0, 1'b0,  8'd13,  9'd173},{  1'b0, 1'b1,  8'd13,  9'd100},
{  1'b0, 1'b0,  8'd87,    9'd0},{  1'b0, 1'b0,  8'd86,    9'd0},{  1'b0, 1'b0,  8'd16,  9'd143},{  1'b0, 1'b1,   8'd0,  9'd176},
{  1'b0, 1'b0,  8'd88,    9'd0},{  1'b0, 1'b0,  8'd87,    9'd0},{  1'b0, 1'b0,  8'd37,    9'd3},{  1'b0, 1'b1,  8'd21,   9'd63},
{  1'b0, 1'b0,  8'd89,    9'd0},{  1'b0, 1'b0,  8'd88,    9'd0},{  1'b0, 1'b0,   8'd9,   9'd28},{  1'b0, 1'b1,   8'd2,   9'd85},
{  1'b0, 1'b0,  8'd90,    9'd0},{  1'b0, 1'b0,  8'd89,    9'd0},{  1'b0, 1'b0,   8'd8,  9'd155},{  1'b0, 1'b1,   8'd5,  9'd136},
{  1'b0, 1'b0,  8'd91,    9'd0},{  1'b0, 1'b0,  8'd90,    9'd0},{  1'b0, 1'b0,  8'd12,  9'd202},{  1'b0, 1'b1,   8'd6,   9'd37},
{  1'b0, 1'b0,  8'd92,    9'd0},{  1'b0, 1'b0,  8'd91,    9'd0},{  1'b0, 1'b0,  8'd19,  9'd359},{  1'b0, 1'b1,   8'd7,  9'd102},
{  1'b0, 1'b0,  8'd93,    9'd0},{  1'b0, 1'b0,  8'd92,    9'd0},{  1'b0, 1'b0,  8'd11,  9'd126},{  1'b0, 1'b1,   8'd6,   9'd76},
{  1'b0, 1'b0,  8'd94,    9'd0},{  1'b0, 1'b0,  8'd93,    9'd0},{  1'b0, 1'b0,  8'd13,  9'd344},{  1'b0, 1'b1,  8'd11,  9'd143},
{  1'b0, 1'b0,  8'd95,    9'd0},{  1'b0, 1'b0,  8'd94,    9'd0},{  1'b0, 1'b0,  8'd31,  9'd166},{  1'b0, 1'b1,   8'd4,  9'd100},
{  1'b0, 1'b0,  8'd96,    9'd0},{  1'b0, 1'b0,  8'd95,    9'd0},{  1'b0, 1'b0,  8'd13,   9'd23},{  1'b0, 1'b1,   8'd7,  9'd278},
{  1'b0, 1'b0,  8'd97,    9'd0},{  1'b0, 1'b0,  8'd96,    9'd0},{  1'b0, 1'b0,   8'd8,   9'd84},{  1'b0, 1'b1,   8'd4,  9'd310},
{  1'b0, 1'b0,  8'd98,    9'd0},{  1'b0, 1'b0,  8'd97,    9'd0},{  1'b0, 1'b0,  8'd13,  9'd262},{  1'b0, 1'b1,   8'd0,  9'd267},
{  1'b0, 1'b0,  8'd99,    9'd0},{  1'b0, 1'b0,  8'd98,    9'd0},{  1'b0, 1'b0,  8'd23,  9'd151},{  1'b0, 1'b1,  8'd11,  9'd112},
{  1'b0, 1'b0, 8'd100,    9'd0},{  1'b0, 1'b0,  8'd99,    9'd0},{  1'b0, 1'b0,  8'd22,  9'd177},{  1'b0, 1'b1,   8'd2,  9'd230},
{  1'b0, 1'b0, 8'd101,    9'd0},{  1'b0, 1'b0, 8'd100,    9'd0},{  1'b0, 1'b0,  8'd37,  9'd200},{  1'b0, 1'b1,  8'd22,  9'd213},
{  1'b0, 1'b0, 8'd102,    9'd0},{  1'b0, 1'b0, 8'd101,    9'd0},{  1'b0, 1'b0,   8'd9,  9'd281},{  1'b0, 1'b1,   8'd6,   9'd65},
{  1'b0, 1'b0, 8'd103,    9'd0},{  1'b0, 1'b0, 8'd102,    9'd0},{  1'b0, 1'b0,  8'd38,  9'd232},{  1'b0, 1'b1,   8'd0,  9'd134},
{  1'b0, 1'b0, 8'd104,    9'd0},{  1'b0, 1'b0, 8'd103,    9'd0},{  1'b0, 1'b0,   8'd3,   9'd45},{  1'b0, 1'b1,   8'd2,  9'd286},
{  1'b0, 1'b0, 8'd105,    9'd0},{  1'b0, 1'b0, 8'd104,    9'd0},{  1'b0, 1'b0,   8'd7,   9'd88},{  1'b0, 1'b1,   8'd0,    9'd8},
{  1'b0, 1'b0, 8'd106,    9'd0},{  1'b0, 1'b0, 8'd105,    9'd0},{  1'b0, 1'b0,  8'd39,   9'd16},{  1'b0, 1'b1,  8'd11,   9'd31},
{  1'b0, 1'b0, 8'd107,    9'd0},{  1'b0, 1'b0, 8'd106,    9'd0},{  1'b0, 1'b0,  8'd15,   9'd61},{  1'b0, 1'b1,   8'd1,  9'd315},
{  1'b0, 1'b0, 8'd108,    9'd0},{  1'b0, 1'b0, 8'd107,    9'd0},{  1'b0, 1'b0,  8'd41,  9'd128},{  1'b0, 1'b1,  8'd14,  9'd317},
{  1'b0, 1'b0, 8'd109,    9'd0},{  1'b0, 1'b0, 8'd108,    9'd0},{  1'b0, 1'b0,  8'd13,   9'd66},{  1'b0, 1'b1,   8'd3,  9'd300},
{  1'b0, 1'b0, 8'd110,    9'd0},{  1'b0, 1'b0, 8'd109,    9'd0},{  1'b0, 1'b0,  8'd11,  9'd319},{  1'b0, 1'b1,   8'd6,  9'd117},
{  1'b0, 1'b0, 8'd111,    9'd0},{  1'b0, 1'b0, 8'd110,    9'd0},{  1'b0, 1'b0,  8'd33,  9'd350},{  1'b0, 1'b1,  8'd13,   9'd43},
{  1'b0, 1'b0, 8'd112,    9'd0},{  1'b0, 1'b0, 8'd111,    9'd0},{  1'b0, 1'b0,  8'd12,  9'd135},{  1'b0, 1'b1,   8'd8,   9'd48},
{  1'b0, 1'b0, 8'd113,    9'd0},{  1'b0, 1'b0, 8'd112,    9'd0},{  1'b0, 1'b0,  8'd38,   9'd89},{  1'b0, 1'b1,  8'd11,   9'd35},
{  1'b0, 1'b0, 8'd114,    9'd0},{  1'b0, 1'b0, 8'd113,    9'd0},{  1'b0, 1'b0,  8'd35,    9'd6},{  1'b0, 1'b1,   8'd9,   9'd42},
{  1'b0, 1'b0, 8'd115,    9'd0},{  1'b0, 1'b0, 8'd114,    9'd0},{  1'b0, 1'b0,  8'd38,  9'd160},{  1'b0, 1'b1,   8'd8,  9'd208},
{  1'b0, 1'b0, 8'd116,    9'd0},{  1'b0, 1'b0, 8'd115,    9'd0},{  1'b0, 1'b0,  8'd26,   9'd52},{  1'b0, 1'b1,   8'd2,  9'd213},
{  1'b0, 1'b0, 8'd117,    9'd0},{  1'b0, 1'b0, 8'd116,    9'd0},{  1'b0, 1'b0,  8'd34,  9'd111},{  1'b0, 1'b1,   8'd4,   9'd59},
{  1'b0, 1'b0, 8'd118,    9'd0},{  1'b0, 1'b0, 8'd117,    9'd0},{  1'b0, 1'b0,   8'd7,   9'd77},{  1'b0, 1'b1,   8'd5,  9'd290},
{  1'b0, 1'b0, 8'd119,    9'd0},{  1'b0, 1'b0, 8'd118,    9'd0},{  1'b0, 1'b0,   8'd4,   9'd98},{  1'b0, 1'b1,   8'd2,  9'd138},
{  1'b0, 1'b0, 8'd120,    9'd0},{  1'b0, 1'b0, 8'd119,    9'd0},{  1'b0, 1'b0,  8'd10,  9'd290},{  1'b0, 1'b1,   8'd9,  9'd201},
{  1'b0, 1'b0, 8'd121,    9'd0},{  1'b0, 1'b0, 8'd120,    9'd0},{  1'b0, 1'b0,  8'd39,  9'd133},{  1'b0, 1'b1,  8'd12,  9'd344},
{  1'b0, 1'b0, 8'd122,    9'd0},{  1'b0, 1'b0, 8'd121,    9'd0},{  1'b0, 1'b0,  8'd12,  9'd219},{  1'b0, 1'b1,   8'd5,   9'd92},
{  1'b0, 1'b0, 8'd123,    9'd0},{  1'b0, 1'b0, 8'd122,    9'd0},{  1'b0, 1'b0,  8'd26,  9'd111},{  1'b0, 1'b1,  8'd14,  9'd285},
{  1'b0, 1'b0, 8'd124,    9'd0},{  1'b0, 1'b0, 8'd123,    9'd0},{  1'b0, 1'b0,  8'd39,    9'd8},{  1'b0, 1'b1,  8'd11,  9'd140},
{  1'b0, 1'b0, 8'd125,    9'd0},{  1'b0, 1'b0, 8'd124,    9'd0},{  1'b0, 1'b0,   8'd6,  9'd338},{  1'b0, 1'b1,   8'd4,  9'd340},
{  1'b0, 1'b0, 8'd126,    9'd0},{  1'b0, 1'b0, 8'd125,    9'd0},{  1'b0, 1'b0,  8'd17,  9'd248},{  1'b0, 1'b1,  8'd11,  9'd218},
{  1'b0, 1'b0, 8'd127,    9'd0},{  1'b0, 1'b0, 8'd126,    9'd0},{  1'b0, 1'b0,  8'd32,   9'd73},{  1'b0, 1'b1,  8'd18,  9'd220},
{  1'b0, 1'b0, 8'd128,    9'd0},{  1'b0, 1'b0, 8'd127,    9'd0},{  1'b0, 1'b0,   8'd5,  9'd329},{  1'b0, 1'b1,   8'd3,  9'd115},
{  1'b0, 1'b0, 8'd129,    9'd0},{  1'b0, 1'b0, 8'd128,    9'd0},{  1'b0, 1'b0,  8'd31,  9'd175},{  1'b0, 1'b1,   8'd1,  9'd121},
{  1'b0, 1'b0, 8'd130,    9'd0},{  1'b0, 1'b0, 8'd129,    9'd0},{  1'b0, 1'b0,  8'd32,  9'd329},{  1'b0, 1'b1,   8'd8,    9'd6},
{  1'b0, 1'b0, 8'd131,    9'd0},{  1'b0, 1'b0, 8'd130,    9'd0},{  1'b0, 1'b0,   8'd8,  9'd190},{  1'b0, 1'b1,   8'd4,  9'd144},
{  1'b0, 1'b0, 8'd132,    9'd0},{  1'b0, 1'b0, 8'd131,    9'd0},{  1'b0, 1'b0,  8'd24,   9'd60},{  1'b0, 1'b1,   8'd7,  9'd243},
{  1'b0, 1'b0, 8'd133,    9'd0},{  1'b0, 1'b0, 8'd132,    9'd0},{  1'b0, 1'b0,   8'd2,  9'd165},{  1'b0, 1'b1,   8'd1,  9'd184},
{  1'b0, 1'b0, 8'd134,    9'd0},{  1'b0, 1'b0, 8'd133,    9'd0},{  1'b0, 1'b0,  8'd12,  9'd123},{  1'b0, 1'b1,   8'd0,  9'd154},
{  1'b0, 1'b0, 8'd135,    9'd0},{  1'b0, 1'b0, 8'd134,    9'd0},{  1'b0, 1'b0,  8'd12,   9'd69},{  1'b0, 1'b1,   8'd8,   9'd49},
{  1'b0, 1'b0, 8'd136,    9'd0},{  1'b0, 1'b0, 8'd135,    9'd0},{  1'b0, 1'b0,  8'd28,   9'd87},{  1'b0, 1'b1,   8'd1,  9'd258},
{  1'b0, 1'b0, 8'd137,    9'd0},{  1'b0, 1'b0, 8'd136,    9'd0},{  1'b0, 1'b0,  8'd37,   9'd34},{  1'b0, 1'b1,  8'd29,  9'd294},
{  1'b0, 1'b0, 8'd138,    9'd0},{  1'b0, 1'b0, 8'd137,    9'd0},{  1'b0, 1'b0,  8'd42,  9'd341},{  1'b0, 1'b1,  8'd18,  9'd218},
{  1'b0, 1'b0, 8'd139,    9'd0},{  1'b0, 1'b0, 8'd138,    9'd0},{  1'b0, 1'b0,  8'd12,  9'd238},{  1'b0, 1'b1,   8'd3,  9'd229},
{  1'b0, 1'b0, 8'd140,    9'd0},{  1'b0, 1'b0, 8'd139,    9'd0},{  1'b0, 1'b0,  8'd41,  9'd181},{  1'b0, 1'b1,  8'd18,  9'd228},
{  1'b0, 1'b0, 8'd141,    9'd0},{  1'b0, 1'b0, 8'd140,    9'd0},{  1'b0, 1'b0,  8'd15,  9'd179},{  1'b0, 1'b1,  8'd12,  9'd262},
{  1'b0, 1'b0, 8'd142,    9'd0},{  1'b0, 1'b0, 8'd141,    9'd0},{  1'b0, 1'b0,  8'd21,  9'd245},{  1'b0, 1'b1,  8'd14,  9'd154},
{  1'b0, 1'b0, 8'd143,    9'd0},{  1'b0, 1'b0, 8'd142,    9'd0},{  1'b0, 1'b0,  8'd19,   9'd68},{  1'b0, 1'b1,   8'd7,  9'd344},
{  1'b0, 1'b0, 8'd144,    9'd0},{  1'b0, 1'b0, 8'd143,    9'd0},{  1'b0, 1'b0,   8'd9,  9'd264},{  1'b0, 1'b1,   8'd2,  9'd103},
{  1'b0, 1'b0, 8'd145,    9'd0},{  1'b0, 1'b0, 8'd144,    9'd0},{  1'b0, 1'b0,  8'd10,   9'd24},{  1'b0, 1'b1,   8'd3,  9'd167},
{  1'b0, 1'b0, 8'd146,    9'd0},{  1'b0, 1'b0, 8'd145,    9'd0},{  1'b0, 1'b0,  8'd31,   9'd82},{  1'b0, 1'b1,   8'd7,   9'd26},
{  1'b0, 1'b0, 8'd147,    9'd0},{  1'b0, 1'b0, 8'd146,    9'd0},{  1'b0, 1'b0,  8'd44,  9'd152},{  1'b0, 1'b1,  8'd13,   9'd53},
{  1'b0, 1'b0, 8'd148,    9'd0},{  1'b0, 1'b0, 8'd147,    9'd0},{  1'b0, 1'b0,  8'd10,  9'd235},{  1'b0, 1'b1,   8'd1,  9'd127},
{  1'b0, 1'b0, 8'd149,    9'd0},{  1'b0, 1'b0, 8'd148,    9'd0},{  1'b0, 1'b0,   8'd5,  9'd295},{  1'b0, 1'b1,   8'd0,  9'd213},
{  1'b0, 1'b0, 8'd150,    9'd0},{  1'b0, 1'b0, 8'd149,    9'd0},{  1'b0, 1'b0,  8'd40,  9'd286},{  1'b0, 1'b1,  8'd27,   9'd40},
{  1'b0, 1'b0, 8'd151,    9'd0},{  1'b0, 1'b0, 8'd150,    9'd0},{  1'b0, 1'b0,  8'd29,  9'd249},{  1'b0, 1'b1,  8'd10,  9'd253},
{  1'b0, 1'b0, 8'd152,    9'd0},{  1'b0, 1'b0, 8'd151,    9'd0},{  1'b0, 1'b0,  8'd14,  9'd305},{  1'b0, 1'b1,  8'd10,   9'd64},
{  1'b0, 1'b0, 8'd153,    9'd0},{  1'b0, 1'b0, 8'd152,    9'd0},{  1'b0, 1'b0,   8'd6,  9'd335},{  1'b0, 1'b1,   8'd0,  9'd348},
{  1'b0, 1'b0, 8'd154,    9'd0},{  1'b0, 1'b0, 8'd153,    9'd0},{  1'b0, 1'b0,  8'd28,  9'd243},{  1'b0, 1'b1,   8'd4,  9'd182},
{  1'b0, 1'b0, 8'd155,    9'd0},{  1'b0, 1'b0, 8'd154,    9'd0},{  1'b0, 1'b0,  8'd44,  9'd345},{  1'b0, 1'b1,  8'd14,  9'd196},
{  1'b0, 1'b0, 8'd156,    9'd0},{  1'b0, 1'b0, 8'd155,    9'd0},{  1'b0, 1'b0,  8'd10,    9'd8},{  1'b0, 1'b1,   8'd6,  9'd143},
{  1'b0, 1'b0, 8'd157,    9'd0},{  1'b0, 1'b0, 8'd156,    9'd0},{  1'b0, 1'b0,  8'd43,  9'd273},{  1'b0, 1'b1,  8'd23,   9'd29},
{  1'b0, 1'b0, 8'd158,    9'd0},{  1'b0, 1'b0, 8'd157,    9'd0},{  1'b0, 1'b0,   8'd9,   9'd51},{  1'b0, 1'b1,   8'd6,  9'd112},
{  1'b0, 1'b0, 8'd159,    9'd0},{  1'b0, 1'b0, 8'd158,    9'd0},{  1'b0, 1'b0,   8'd3,  9'd164},{  1'b0, 1'b1,   8'd3,  9'd124},
{  1'b0, 1'b0, 8'd160,    9'd0},{  1'b0, 1'b0, 8'd159,    9'd0},{  1'b0, 1'b0,  8'd20,   9'd30},{  1'b0, 1'b1,   8'd9,   9'd80},
{  1'b0, 1'b0, 8'd161,    9'd0},{  1'b0, 1'b0, 8'd160,    9'd0},{  1'b0, 1'b0,  8'd32,  9'd255},{  1'b0, 1'b1,   8'd0,  9'd174},
{  1'b0, 1'b0, 8'd162,    9'd0},{  1'b0, 1'b0, 8'd161,    9'd0},{  1'b0, 1'b0,  8'd13,  9'd115},{  1'b0, 1'b1,   8'd1,  9'd155},
{  1'b0, 1'b0, 8'd163,    9'd0},{  1'b0, 1'b0, 8'd162,    9'd0},{  1'b0, 1'b0,  8'd10,   9'd93},{  1'b0, 1'b1,   8'd1,  9'd124},
{  1'b0, 1'b0, 8'd164,    9'd0},{  1'b0, 1'b0, 8'd163,    9'd0},{  1'b0, 1'b0,  8'd14,   9'd10},{  1'b0, 1'b1,   8'd2,   9'd13},
{  1'b0, 1'b0, 8'd165,    9'd0},{  1'b0, 1'b0, 8'd164,    9'd0},{  1'b0, 1'b0,  8'd43,  9'd135},{  1'b0, 1'b1,  8'd21,  9'd254},
{  1'b0, 1'b0, 8'd166,    9'd0},{  1'b0, 1'b0, 8'd165,    9'd0},{  1'b0, 1'b0,  8'd26,  9'd337},{  1'b0, 1'b1,  8'd10,  9'd123},
{  1'b0, 1'b0, 8'd167,    9'd0},{  1'b0, 1'b0, 8'd166,    9'd0},{  1'b0, 1'b0,  8'd34,  9'd336},{  1'b0, 1'b1,   8'd3,  9'd166},
{  1'b0, 1'b0, 8'd168,    9'd0},{  1'b0, 1'b0, 8'd167,    9'd0},{  1'b0, 1'b0,  8'd43,  9'd150},{  1'b0, 1'b1,  8'd16,   9'd73},
{  1'b0, 1'b0, 8'd169,    9'd0},{  1'b0, 1'b0, 8'd168,    9'd0},{  1'b0, 1'b0,  8'd42,  9'd229},{  1'b0, 1'b1,   8'd7,  9'd238},
{  1'b0, 1'b0, 8'd170,    9'd0},{  1'b0, 1'b0, 8'd169,    9'd0},{  1'b0, 1'b0,  8'd22,  9'd166},{  1'b0, 1'b1,  8'd14,  9'd201},
{  1'b0, 1'b0, 8'd171,    9'd0},{  1'b0, 1'b0, 8'd170,    9'd0},{  1'b0, 1'b0,  8'd20,  9'd281},{  1'b0, 1'b1,   8'd4,  9'd242},
{  1'b0, 1'b0, 8'd172,    9'd0},{  1'b0, 1'b0, 8'd171,    9'd0},{  1'b0, 1'b0,  8'd30,  9'd221},{  1'b0, 1'b1,  8'd16,  9'd205},
{  1'b0, 1'b0, 8'd173,    9'd0},{  1'b0, 1'b0, 8'd172,    9'd0},{  1'b0, 1'b0,  8'd13,  9'd197},{  1'b0, 1'b1,   8'd5,  9'd257},
{  1'b0, 1'b0, 8'd174,    9'd0},{  1'b0, 1'b0, 8'd173,    9'd0},{  1'b0, 1'b0,  8'd25,  9'd158},{  1'b0, 1'b1,  8'd14,  9'd347},
{  1'b0, 1'b0, 8'd175,    9'd0},{  1'b0, 1'b0, 8'd174,    9'd0},{  1'b0, 1'b0,  8'd33,  9'd103},{  1'b0, 1'b1,   8'd7,   9'd10},
{  1'b0, 1'b0, 8'd176,    9'd0},{  1'b0, 1'b0, 8'd175,    9'd0},{  1'b0, 1'b0,   8'd5,   9'd72},{  1'b0, 1'b1,   8'd3,   9'd67},
{  1'b0, 1'b0, 8'd177,    9'd0},{  1'b0, 1'b0, 8'd176,    9'd0},{  1'b0, 1'b0,   8'd9,  9'd162},{  1'b0, 1'b1,   8'd3,  9'd176},
{  1'b0, 1'b0, 8'd178,    9'd0},{  1'b0, 1'b0, 8'd177,    9'd0},{  1'b0, 1'b0,   8'd7,   9'd50},{  1'b0, 1'b1,   8'd1,   9'd56},
{  1'b0, 1'b0, 8'd179,    9'd0},{  1'b0, 1'b0, 8'd178,    9'd0},{  1'b0, 1'b0,  8'd36,   9'd98},{  1'b0, 1'b1,   8'd2,  9'd296}
};
localparam bit [18 : 0] cLARGE_HS_V_TAB_1BY4_PACKED[cLARGE_HS_TAB_1BY4_PACKED_SIZE] = '{
{8'd179, 1'b0,   10'd0},{8'd179, 1'b1, 10'd536},
{8'd178, 1'b0, 10'd532},{8'd178, 1'b1, 10'd537},
{8'd177, 1'b0, 10'd528},{8'd177, 1'b1, 10'd533},
{8'd176, 1'b0, 10'd524},{8'd176, 1'b1, 10'd529},
{8'd175, 1'b0, 10'd520},{8'd175, 1'b1, 10'd525},
{8'd174, 1'b0, 10'd516},{8'd174, 1'b1, 10'd521},
{8'd173, 1'b0, 10'd512},{8'd173, 1'b1, 10'd517},
{8'd172, 1'b0, 10'd508},{8'd172, 1'b1, 10'd513},
{8'd171, 1'b0, 10'd504},{8'd171, 1'b1, 10'd509},
{8'd170, 1'b0, 10'd500},{8'd170, 1'b1, 10'd505},
{8'd169, 1'b0, 10'd496},{8'd169, 1'b1, 10'd501},
{8'd168, 1'b0, 10'd492},{8'd168, 1'b1, 10'd497},
{8'd167, 1'b0, 10'd488},{8'd167, 1'b1, 10'd493},
{8'd166, 1'b0, 10'd484},{8'd166, 1'b1, 10'd489},
{8'd165, 1'b0, 10'd480},{8'd165, 1'b1, 10'd485},
{8'd164, 1'b0, 10'd476},{8'd164, 1'b1, 10'd481},
{8'd163, 1'b0, 10'd472},{8'd163, 1'b1, 10'd477},
{8'd162, 1'b0, 10'd468},{8'd162, 1'b1, 10'd473},
{8'd161, 1'b0, 10'd464},{8'd161, 1'b1, 10'd469},
{8'd160, 1'b0, 10'd460},{8'd160, 1'b1, 10'd465},
{8'd159, 1'b0, 10'd456},{8'd159, 1'b1, 10'd461},
{8'd158, 1'b0, 10'd452},{8'd158, 1'b1, 10'd457},
{8'd157, 1'b0, 10'd448},{8'd157, 1'b1, 10'd453},
{8'd156, 1'b0, 10'd444},{8'd156, 1'b1, 10'd449},
{8'd155, 1'b0, 10'd440},{8'd155, 1'b1, 10'd445},
{8'd154, 1'b0, 10'd436},{8'd154, 1'b1, 10'd441},
{8'd153, 1'b0, 10'd432},{8'd153, 1'b1, 10'd437},
{8'd152, 1'b0, 10'd428},{8'd152, 1'b1, 10'd433},
{8'd151, 1'b0, 10'd424},{8'd151, 1'b1, 10'd429},
{8'd150, 1'b0, 10'd420},{8'd150, 1'b1, 10'd425},
{8'd149, 1'b0, 10'd416},{8'd149, 1'b1, 10'd421},
{8'd148, 1'b0, 10'd412},{8'd148, 1'b1, 10'd417},
{8'd147, 1'b0, 10'd408},{8'd147, 1'b1, 10'd413},
{8'd146, 1'b0, 10'd404},{8'd146, 1'b1, 10'd409},
{8'd145, 1'b0, 10'd400},{8'd145, 1'b1, 10'd405},
{8'd144, 1'b0, 10'd396},{8'd144, 1'b1, 10'd401},
{8'd143, 1'b0, 10'd392},{8'd143, 1'b1, 10'd397},
{8'd142, 1'b0, 10'd388},{8'd142, 1'b1, 10'd393},
{8'd141, 1'b0, 10'd384},{8'd141, 1'b1, 10'd389},
{8'd140, 1'b0, 10'd380},{8'd140, 1'b1, 10'd385},
{8'd139, 1'b0, 10'd376},{8'd139, 1'b1, 10'd381},
{8'd138, 1'b0, 10'd372},{8'd138, 1'b1, 10'd377},
{8'd137, 1'b0, 10'd368},{8'd137, 1'b1, 10'd373},
{8'd136, 1'b0, 10'd364},{8'd136, 1'b1, 10'd369},
{8'd135, 1'b0, 10'd360},{8'd135, 1'b1, 10'd365},
{8'd134, 1'b0, 10'd356},{8'd134, 1'b1, 10'd361},
{8'd133, 1'b0, 10'd352},{8'd133, 1'b1, 10'd357},
{8'd132, 1'b0, 10'd348},{8'd132, 1'b1, 10'd353},
{8'd131, 1'b0, 10'd344},{8'd131, 1'b1, 10'd349},
{8'd130, 1'b0, 10'd340},{8'd130, 1'b1, 10'd345},
{8'd129, 1'b0, 10'd336},{8'd129, 1'b1, 10'd341},
{8'd128, 1'b0, 10'd332},{8'd128, 1'b1, 10'd337},
{8'd127, 1'b0, 10'd328},{8'd127, 1'b1, 10'd333},
{8'd126, 1'b0, 10'd324},{8'd126, 1'b1, 10'd329},
{8'd125, 1'b0, 10'd320},{8'd125, 1'b1, 10'd325},
{8'd124, 1'b0, 10'd316},{8'd124, 1'b1, 10'd321},
{8'd123, 1'b0, 10'd312},{8'd123, 1'b1, 10'd317},
{8'd122, 1'b0, 10'd308},{8'd122, 1'b1, 10'd313},
{8'd121, 1'b0, 10'd304},{8'd121, 1'b1, 10'd309},
{8'd120, 1'b0, 10'd300},{8'd120, 1'b1, 10'd305},
{8'd119, 1'b0, 10'd296},{8'd119, 1'b1, 10'd301},
{8'd118, 1'b0, 10'd292},{8'd118, 1'b1, 10'd297},
{8'd117, 1'b0, 10'd288},{8'd117, 1'b1, 10'd293},
{8'd116, 1'b0, 10'd284},{8'd116, 1'b1, 10'd289},
{8'd115, 1'b0, 10'd280},{8'd115, 1'b1, 10'd285},
{8'd114, 1'b0, 10'd276},{8'd114, 1'b1, 10'd281},
{8'd113, 1'b0, 10'd272},{8'd113, 1'b1, 10'd277},
{8'd112, 1'b0, 10'd268},{8'd112, 1'b1, 10'd273},
{8'd111, 1'b0, 10'd264},{8'd111, 1'b1, 10'd269},
{8'd110, 1'b0, 10'd260},{8'd110, 1'b1, 10'd265},
{8'd109, 1'b0, 10'd256},{8'd109, 1'b1, 10'd261},
{8'd108, 1'b0, 10'd252},{8'd108, 1'b1, 10'd257},
{8'd107, 1'b0, 10'd248},{8'd107, 1'b1, 10'd253},
{8'd106, 1'b0, 10'd244},{8'd106, 1'b1, 10'd249},
{8'd105, 1'b0, 10'd240},{8'd105, 1'b1, 10'd245},
{8'd104, 1'b0, 10'd236},{8'd104, 1'b1, 10'd241},
{8'd103, 1'b0, 10'd232},{8'd103, 1'b1, 10'd237},
{8'd102, 1'b0, 10'd228},{8'd102, 1'b1, 10'd233},
{8'd101, 1'b0, 10'd224},{8'd101, 1'b1, 10'd229},
{8'd100, 1'b0, 10'd220},{8'd100, 1'b1, 10'd225},
{ 8'd99, 1'b0, 10'd216},{ 8'd99, 1'b1, 10'd221},
{ 8'd98, 1'b0, 10'd212},{ 8'd98, 1'b1, 10'd217},
{ 8'd97, 1'b0, 10'd208},{ 8'd97, 1'b1, 10'd213},
{ 8'd96, 1'b0, 10'd204},{ 8'd96, 1'b1, 10'd209},
{ 8'd95, 1'b0, 10'd200},{ 8'd95, 1'b1, 10'd205},
{ 8'd94, 1'b0, 10'd196},{ 8'd94, 1'b1, 10'd201},
{ 8'd93, 1'b0, 10'd192},{ 8'd93, 1'b1, 10'd197},
{ 8'd92, 1'b0, 10'd188},{ 8'd92, 1'b1, 10'd193},
{ 8'd91, 1'b0, 10'd184},{ 8'd91, 1'b1, 10'd189},
{ 8'd90, 1'b0, 10'd180},{ 8'd90, 1'b1, 10'd185},
{ 8'd89, 1'b0, 10'd176},{ 8'd89, 1'b1, 10'd181},
{ 8'd88, 1'b0, 10'd172},{ 8'd88, 1'b1, 10'd177},
{ 8'd87, 1'b0, 10'd168},{ 8'd87, 1'b1, 10'd173},
{ 8'd86, 1'b0, 10'd164},{ 8'd86, 1'b1, 10'd169},
{ 8'd85, 1'b0, 10'd160},{ 8'd85, 1'b1, 10'd165},
{ 8'd84, 1'b0, 10'd156},{ 8'd84, 1'b1, 10'd161},
{ 8'd83, 1'b0, 10'd152},{ 8'd83, 1'b1, 10'd157},
{ 8'd82, 1'b0, 10'd148},{ 8'd82, 1'b1, 10'd153},
{ 8'd81, 1'b0, 10'd144},{ 8'd81, 1'b1, 10'd149},
{ 8'd80, 1'b0, 10'd140},{ 8'd80, 1'b1, 10'd145},
{ 8'd79, 1'b0, 10'd136},{ 8'd79, 1'b1, 10'd141},
{ 8'd78, 1'b0, 10'd132},{ 8'd78, 1'b1, 10'd137},
{ 8'd77, 1'b0, 10'd128},{ 8'd77, 1'b1, 10'd133},
{ 8'd76, 1'b0, 10'd124},{ 8'd76, 1'b1, 10'd129},
{ 8'd75, 1'b0, 10'd120},{ 8'd75, 1'b1, 10'd125},
{ 8'd74, 1'b0, 10'd116},{ 8'd74, 1'b1, 10'd121},
{ 8'd73, 1'b0, 10'd112},{ 8'd73, 1'b1, 10'd117},
{ 8'd72, 1'b0, 10'd108},{ 8'd72, 1'b1, 10'd113},
{ 8'd71, 1'b0, 10'd104},{ 8'd71, 1'b1, 10'd109},
{ 8'd70, 1'b0, 10'd100},{ 8'd70, 1'b1, 10'd105},
{ 8'd69, 1'b0,  10'd96},{ 8'd69, 1'b1, 10'd101},
{ 8'd68, 1'b0,  10'd92},{ 8'd68, 1'b1,  10'd97},
{ 8'd67, 1'b0,  10'd88},{ 8'd67, 1'b1,  10'd93},
{ 8'd66, 1'b0,  10'd84},{ 8'd66, 1'b1,  10'd89},
{ 8'd65, 1'b0,  10'd80},{ 8'd65, 1'b1,  10'd85},
{ 8'd64, 1'b0,  10'd76},{ 8'd64, 1'b1,  10'd81},
{ 8'd63, 1'b0,  10'd72},{ 8'd63, 1'b1,  10'd77},
{ 8'd62, 1'b0,  10'd68},{ 8'd62, 1'b1,  10'd73},
{ 8'd61, 1'b0,  10'd64},{ 8'd61, 1'b1,  10'd69},
{ 8'd60, 1'b0,  10'd60},{ 8'd60, 1'b1,  10'd65},
{ 8'd59, 1'b0,  10'd56},{ 8'd59, 1'b1,  10'd61},
{ 8'd58, 1'b0,  10'd52},{ 8'd58, 1'b1,  10'd57},
{ 8'd57, 1'b0,  10'd48},{ 8'd57, 1'b1,  10'd53},
{ 8'd56, 1'b0,  10'd44},{ 8'd56, 1'b1,  10'd49},
{ 8'd55, 1'b0,  10'd40},{ 8'd55, 1'b1,  10'd45},
{ 8'd54, 1'b0,  10'd36},{ 8'd54, 1'b1,  10'd41},
{ 8'd53, 1'b0,  10'd32},{ 8'd53, 1'b1,  10'd37},
{ 8'd52, 1'b0,  10'd28},{ 8'd52, 1'b1,  10'd33},
{ 8'd51, 1'b0,  10'd24},{ 8'd51, 1'b1,  10'd29},
{ 8'd50, 1'b0,  10'd20},{ 8'd50, 1'b1,  10'd25},
{ 8'd49, 1'b0,  10'd16},{ 8'd49, 1'b1,  10'd21},
{ 8'd48, 1'b0,  10'd12},{ 8'd48, 1'b1,  10'd17},
{ 8'd47, 1'b0,   10'd8},{ 8'd47, 1'b1,  10'd13},
{ 8'd46, 1'b0,   10'd4},{ 8'd46, 1'b1,   10'd9},
{ 8'd45, 1'b0,   10'd1},{ 8'd45, 1'b1,   10'd5},
{ 8'd44, 1'b0,   10'd6},{ 8'd44, 1'b0, 10'd410},{ 8'd44, 1'b1, 10'd442},
{ 8'd43, 1'b0, 10'd450},{ 8'd43, 1'b0, 10'd482},{ 8'd43, 1'b1, 10'd494},
{ 8'd42, 1'b0,  10'd54},{ 8'd42, 1'b0, 10'd374},{ 8'd42, 1'b1, 10'd498},
{ 8'd41, 1'b0,  10'd38},{ 8'd41, 1'b0, 10'd254},{ 8'd41, 1'b1, 10'd382},
{ 8'd40, 1'b0,  10'd74},{ 8'd40, 1'b0, 10'd142},{ 8'd40, 1'b1, 10'd422},
{ 8'd39, 1'b0, 10'd246},{ 8'd39, 1'b0, 10'd306},{ 8'd39, 1'b1, 10'd318},
{ 8'd38, 1'b0, 10'd234},{ 8'd38, 1'b0, 10'd274},{ 8'd38, 1'b1, 10'd282},
{ 8'd37, 1'b0, 10'd174},{ 8'd37, 1'b0, 10'd226},{ 8'd37, 1'b1, 10'd370},
{ 8'd36, 1'b0,  10'd94},{ 8'd36, 1'b0, 10'd130},{ 8'd36, 1'b1, 10'd538},
{ 8'd35, 1'b0,  10'd34},{ 8'd35, 1'b0,  10'd90},{ 8'd35, 1'b1, 10'd278},
{ 8'd34, 1'b0, 10'd106},{ 8'd34, 1'b0, 10'd290},{ 8'd34, 1'b1, 10'd490},
{ 8'd33, 1'b0, 10'd162},{ 8'd33, 1'b0, 10'd266},{ 8'd33, 1'b1, 10'd522},
{ 8'd32, 1'b0, 10'd330},{ 8'd32, 1'b0, 10'd342},{ 8'd32, 1'b1, 10'd466},
{ 8'd31, 1'b0, 10'd202},{ 8'd31, 1'b0, 10'd338},{ 8'd31, 1'b1, 10'd406},
{ 8'd30, 1'b0,  10'd82},{ 8'd30, 1'b0, 10'd122},{ 8'd30, 1'b1, 10'd510},
{ 8'd29, 1'b0,  10'd58},{ 8'd29, 1'b0, 10'd371},{ 8'd29, 1'b1, 10'd426},
{ 8'd28, 1'b0,   10'd7},{ 8'd28, 1'b0, 10'd366},{ 8'd28, 1'b1, 10'd438},
{ 8'd27, 1'b0,   10'd2},{ 8'd27, 1'b0, 10'd154},{ 8'd27, 1'b1, 10'd423},
{ 8'd26, 1'b0, 10'd286},{ 8'd26, 1'b0, 10'd314},{ 8'd26, 1'b1, 10'd486},
{ 8'd25, 1'b0,  10'd22},{ 8'd25, 1'b0, 10'd134},{ 8'd25, 1'b1, 10'd518},
{ 8'd24, 1'b0,  10'd35},{ 8'd24, 1'b0, 10'd131},{ 8'd24, 1'b1, 10'd350},
{ 8'd23, 1'b0,  10'd86},{ 8'd23, 1'b0, 10'd218},{ 8'd23, 1'b1, 10'd451},
{ 8'd22, 1'b0, 10'd222},{ 8'd22, 1'b0, 10'd227},{ 8'd22, 1'b1, 10'd502},
{ 8'd21, 1'b0, 10'd175},{ 8'd21, 1'b0, 10'd390},{ 8'd21, 1'b1, 10'd483},
{ 8'd20, 1'b0,  10'd14},{ 8'd20, 1'b0, 10'd462},{ 8'd20, 1'b1, 10'd506},
{ 8'd19, 1'b0, 10'd158},{ 8'd19, 1'b0, 10'd190},{ 8'd19, 1'b1, 10'd394},
{ 8'd18, 1'b0, 10'd331},{ 8'd18, 1'b0, 10'd375},{ 8'd18, 1'b1, 10'd383},
{ 8'd17, 1'b0,  10'd39},{ 8'd17, 1'b0, 10'd107},{ 8'd17, 1'b1, 10'd326},
{ 8'd16, 1'b0, 10'd170},{ 8'd16, 1'b0, 10'd495},{ 8'd16, 1'b1, 10'd511},
{ 8'd15, 1'b0,  10'd50},{ 8'd15, 1'b0, 10'd250},{ 8'd15, 1'b1, 10'd386},
{ 8'd14, 1'b0,  10'd10},{ 8'd14, 1'b0,  10'd55},{ 8'd14, 1'b0,  10'd87},{ 8'd14, 1'b0, 10'd114},{ 8'd14, 1'b0, 10'd255},{ 8'd14, 1'b0, 10'd315},{ 8'd14, 1'b0, 10'd391},{ 8'd14, 1'b0, 10'd430},{ 8'd14, 1'b0, 10'd443},{ 8'd14, 1'b0, 10'd478},{ 8'd14, 1'b0, 10'd503},{ 8'd14, 1'b1, 10'd519},
{ 8'd13, 1'b0,  10'd15},{ 8'd13, 1'b0, 10'd102},{ 8'd13, 1'b0, 10'd166},{ 8'd13, 1'b0, 10'd167},{ 8'd13, 1'b0, 10'd198},{ 8'd13, 1'b0, 10'd206},{ 8'd13, 1'b0, 10'd214},{ 8'd13, 1'b0, 10'd258},{ 8'd13, 1'b0, 10'd267},{ 8'd13, 1'b0, 10'd411},{ 8'd13, 1'b0, 10'd470},{ 8'd13, 1'b1, 10'd514},
{ 8'd12, 1'b0,  10'd30},{ 8'd12, 1'b0,  10'd46},{ 8'd12, 1'b0,  10'd70},{ 8'd12, 1'b0,  10'd78},{ 8'd12, 1'b0, 10'd186},{ 8'd12, 1'b0, 10'd270},{ 8'd12, 1'b0, 10'd307},{ 8'd12, 1'b0, 10'd310},{ 8'd12, 1'b0, 10'd358},{ 8'd12, 1'b0, 10'd362},{ 8'd12, 1'b0, 10'd378},{ 8'd12, 1'b1, 10'd387},
{ 8'd11, 1'b0,  10'd18},{ 8'd11, 1'b0,  10'd59},{ 8'd11, 1'b0,  10'd83},{ 8'd11, 1'b0, 10'd135},{ 8'd11, 1'b0, 10'd194},{ 8'd11, 1'b0, 10'd199},{ 8'd11, 1'b0, 10'd219},{ 8'd11, 1'b0, 10'd247},{ 8'd11, 1'b0, 10'd262},{ 8'd11, 1'b0, 10'd275},{ 8'd11, 1'b0, 10'd319},{ 8'd11, 1'b1, 10'd327},
{ 8'd10, 1'b0,  10'd31},{ 8'd10, 1'b0,  10'd42},{ 8'd10, 1'b0,  10'd95},{ 8'd10, 1'b0, 10'd143},{ 8'd10, 1'b0, 10'd302},{ 8'd10, 1'b0, 10'd402},{ 8'd10, 1'b0, 10'd414},{ 8'd10, 1'b0, 10'd427},{ 8'd10, 1'b0, 10'd431},{ 8'd10, 1'b0, 10'd446},{ 8'd10, 1'b0, 10'd474},{ 8'd10, 1'b1, 10'd487},
{  8'd9, 1'b0,  10'd43},{  8'd9, 1'b0,  10'd75},{  8'd9, 1'b0, 10'd150},{  8'd9, 1'b0, 10'd159},{  8'd9, 1'b0, 10'd178},{  8'd9, 1'b0, 10'd230},{  8'd9, 1'b0, 10'd279},{  8'd9, 1'b0, 10'd303},{  8'd9, 1'b0, 10'd398},{  8'd9, 1'b0, 10'd454},{  8'd9, 1'b0, 10'd463},{  8'd9, 1'b1, 10'd530},
{  8'd8, 1'b0,  10'd51},{  8'd8, 1'b0,  10'd71},{  8'd8, 1'b0,  10'd79},{  8'd8, 1'b0,  10'd98},{  8'd8, 1'b0, 10'd138},{  8'd8, 1'b0, 10'd182},{  8'd8, 1'b0, 10'd210},{  8'd8, 1'b0, 10'd271},{  8'd8, 1'b0, 10'd283},{  8'd8, 1'b0, 10'd343},{  8'd8, 1'b0, 10'd346},{  8'd8, 1'b1, 10'd363},
{  8'd7, 1'b0,  10'd66},{  8'd7, 1'b0, 10'd115},{  8'd7, 1'b0, 10'd191},{  8'd7, 1'b0, 10'd207},{  8'd7, 1'b0, 10'd242},{  8'd7, 1'b0, 10'd294},{  8'd7, 1'b0, 10'd351},{  8'd7, 1'b0, 10'd395},{  8'd7, 1'b0, 10'd407},{  8'd7, 1'b0, 10'd499},{  8'd7, 1'b0, 10'd523},{  8'd7, 1'b1, 10'd534},
{  8'd6, 1'b0,  10'd11},{  8'd6, 1'b0,  10'd99},{  8'd6, 1'b0, 10'd123},{  8'd6, 1'b0, 10'd146},{  8'd6, 1'b0, 10'd187},{  8'd6, 1'b0, 10'd195},{  8'd6, 1'b0, 10'd231},{  8'd6, 1'b0, 10'd263},{  8'd6, 1'b0, 10'd322},{  8'd6, 1'b0, 10'd434},{  8'd6, 1'b0, 10'd447},{  8'd6, 1'b1, 10'd455},
{  8'd5, 1'b0,  10'd26},{  8'd5, 1'b0,  10'd27},{  8'd5, 1'b0, 10'd103},{  8'd5, 1'b0, 10'd126},{  8'd5, 1'b0, 10'd163},{  8'd5, 1'b0, 10'd183},{  8'd5, 1'b0, 10'd295},{  8'd5, 1'b0, 10'd311},{  8'd5, 1'b0, 10'd334},{  8'd5, 1'b0, 10'd418},{  8'd5, 1'b0, 10'd515},{  8'd5, 1'b1, 10'd526},
{  8'd4, 1'b0,  10'd23},{  8'd4, 1'b0, 10'd110},{  8'd4, 1'b0, 10'd127},{  8'd4, 1'b0, 10'd147},{  8'd4, 1'b0, 10'd203},{  8'd4, 1'b0, 10'd211},{  8'd4, 1'b0, 10'd291},{  8'd4, 1'b0, 10'd298},{  8'd4, 1'b0, 10'd323},{  8'd4, 1'b0, 10'd347},{  8'd4, 1'b0, 10'd439},{  8'd4, 1'b1, 10'd507},
{  8'd3, 1'b0, 10'd111},{  8'd3, 1'b0, 10'd155},{  8'd3, 1'b0, 10'd238},{  8'd3, 1'b0, 10'd259},{  8'd3, 1'b0, 10'd335},{  8'd3, 1'b0, 10'd379},{  8'd3, 1'b0, 10'd403},{  8'd3, 1'b0, 10'd458},{  8'd3, 1'b0, 10'd459},{  8'd3, 1'b0, 10'd491},{  8'd3, 1'b0, 10'd527},{  8'd3, 1'b1, 10'd531},
{  8'd2, 1'b0,  10'd47},{  8'd2, 1'b0,  10'd62},{  8'd2, 1'b0, 10'd118},{  8'd2, 1'b0, 10'd179},{  8'd2, 1'b0, 10'd223},{  8'd2, 1'b0, 10'd239},{  8'd2, 1'b0, 10'd287},{  8'd2, 1'b0, 10'd299},{  8'd2, 1'b0, 10'd354},{  8'd2, 1'b0, 10'd399},{  8'd2, 1'b0, 10'd479},{  8'd2, 1'b1, 10'd539},
{  8'd1, 1'b0,  10'd19},{  8'd1, 1'b0,  10'd91},{  8'd1, 1'b0, 10'd139},{  8'd1, 1'b0, 10'd151},{  8'd1, 1'b0, 10'd251},{  8'd1, 1'b0, 10'd339},{  8'd1, 1'b0, 10'd355},{  8'd1, 1'b0, 10'd367},{  8'd1, 1'b0, 10'd415},{  8'd1, 1'b0, 10'd471},{  8'd1, 1'b0, 10'd475},{  8'd1, 1'b1, 10'd535},
{  8'd0, 1'b0,   10'd3},{  8'd0, 1'b0,  10'd63},{  8'd0, 1'b0,  10'd67},{  8'd0, 1'b0, 10'd119},{  8'd0, 1'b0, 10'd171},{  8'd0, 1'b0, 10'd215},{  8'd0, 1'b0, 10'd235},{  8'd0, 1'b0, 10'd243},{  8'd0, 1'b0, 10'd359},{  8'd0, 1'b0, 10'd419},{  8'd0, 1'b0, 10'd435},{  8'd0, 1'b1, 10'd467}
};
localparam int          cLARGE_HS_TAB_1BY3_PACKED_SIZE = 600;
localparam bit [18 : 0] cLARGE_HS_TAB_1BY3_PACKED[cLARGE_HS_TAB_1BY3_PACKED_SIZE] = '{
{  1'b1, 1'b0, 8'd179,    9'd1},{  1'b0, 1'b0,  8'd60,    9'd0},{  1'b0, 1'b0,  8'd44,  9'd313},{  1'b0, 1'b0,   8'd0,   9'd46},{  1'b0, 1'b1,   8'd0,  9'd176},
{  1'b0, 1'b0,  8'd61,    9'd0},{  1'b0, 1'b0,  8'd60,    9'd0},{  1'b0, 1'b0,  8'd54,  9'd236},{  1'b0, 1'b0,  8'd46,  9'd184},{  1'b0, 1'b1,  8'd35,  9'd228},
{  1'b0, 1'b0,  8'd62,    9'd0},{  1'b0, 1'b0,  8'd61,    9'd0},{  1'b0, 1'b0,  8'd27,  9'd284},{  1'b0, 1'b0,  8'd16,  9'd243},{  1'b0, 1'b1,   8'd6,  9'd143},
{  1'b0, 1'b0,  8'd63,    9'd0},{  1'b0, 1'b0,  8'd62,    9'd0},{  1'b0, 1'b0,  8'd46,  9'd209},{  1'b0, 1'b0,  8'd12,  9'd332},{  1'b0, 1'b1,   8'd1,  9'd123},
{  1'b0, 1'b0,  8'd64,    9'd0},{  1'b0, 1'b0,  8'd63,    9'd0},{  1'b0, 1'b0,  8'd23,  9'd345},{  1'b0, 1'b0,  8'd13,   9'd20},{  1'b0, 1'b1,  8'd10,  9'd355},
{  1'b0, 1'b0,  8'd65,    9'd0},{  1'b0, 1'b0,  8'd64,    9'd0},{  1'b0, 1'b0,  8'd18,   9'd16},{  1'b0, 1'b0,  8'd17,   9'd86},{  1'b0, 1'b1,   8'd4,  9'd201},
{  1'b0, 1'b0,  8'd66,    9'd0},{  1'b0, 1'b0,  8'd65,    9'd0},{  1'b0, 1'b0,  8'd15,  9'd263},{  1'b0, 1'b0,   8'd5,  9'd103},{  1'b0, 1'b1,   8'd5,  9'd189},
{  1'b0, 1'b0,  8'd67,    9'd0},{  1'b0, 1'b0,  8'd66,    9'd0},{  1'b0, 1'b0,  8'd47,   9'd67},{  1'b0, 1'b0,  8'd18,  9'd128},{  1'b0, 1'b1,   8'd9,  9'd101},
{  1'b0, 1'b0,  8'd68,    9'd0},{  1'b0, 1'b0,  8'd67,    9'd0},{  1'b0, 1'b0,  8'd34,  9'd330},{  1'b0, 1'b0,  8'd22,  9'd133},{  1'b0, 1'b1,  8'd21,  9'd145},
{  1'b0, 1'b0,  8'd69,    9'd0},{  1'b0, 1'b0,  8'd68,    9'd0},{  1'b0, 1'b0,  8'd23,  9'd227},{  1'b0, 1'b0,  8'd16,   9'd54},{  1'b0, 1'b1,   8'd9,  9'd289},
{  1'b0, 1'b0,  8'd70,    9'd0},{  1'b0, 1'b0,  8'd69,    9'd0},{  1'b0, 1'b0,  8'd45,  9'd263},{  1'b0, 1'b0,  8'd19,  9'd177},{  1'b0, 1'b1,   8'd2,   9'd97},
{  1'b0, 1'b0,  8'd71,    9'd0},{  1'b0, 1'b0,  8'd70,    9'd0},{  1'b0, 1'b0,  8'd16,  9'd108},{  1'b0, 1'b0,   8'd9,   9'd63},{  1'b0, 1'b1,   8'd8,  9'd312},
{  1'b0, 1'b0,  8'd72,    9'd0},{  1'b0, 1'b0,  8'd71,    9'd0},{  1'b0, 1'b0,  8'd54,   9'd41},{  1'b0, 1'b0,  8'd16,  9'd311},{  1'b0, 1'b1,  8'd14,  9'd151},
{  1'b0, 1'b0,  8'd73,    9'd0},{  1'b0, 1'b0,  8'd72,    9'd0},{  1'b0, 1'b0,  8'd11,   9'd62},{  1'b0, 1'b0,  8'd10,  9'd144},{  1'b0, 1'b1,   8'd0,  9'd134},
{  1'b0, 1'b0,  8'd74,    9'd0},{  1'b0, 1'b0,  8'd73,    9'd0},{  1'b0, 1'b0,  8'd22,  9'd323},{  1'b0, 1'b0,   8'd2,  9'd224},{  1'b0, 1'b1,   8'd0,  9'd137},
{  1'b0, 1'b0,  8'd75,    9'd0},{  1'b0, 1'b0,  8'd74,    9'd0},{  1'b0, 1'b0,  8'd44,  9'd119},{  1'b0, 1'b0,  8'd11,   9'd92},{  1'b0, 1'b1,   8'd7,  9'd328},
{  1'b0, 1'b0,  8'd76,    9'd0},{  1'b0, 1'b0,  8'd75,    9'd0},{  1'b0, 1'b0,  8'd57,   9'd66},{  1'b0, 1'b0,  8'd52,   9'd10},{  1'b0, 1'b1,  8'd17,    9'd6},
{  1'b0, 1'b0,  8'd77,    9'd0},{  1'b0, 1'b0,  8'd76,    9'd0},{  1'b0, 1'b0,  8'd35,  9'd245},{  1'b0, 1'b0,  8'd34,  9'd176},{  1'b0, 1'b1,  8'd13,  9'd237},
{  1'b0, 1'b0,  8'd78,    9'd0},{  1'b0, 1'b0,  8'd77,    9'd0},{  1'b0, 1'b0,  8'd58,   9'd88},{  1'b0, 1'b0,   8'd8,  9'd206},{  1'b0, 1'b1,   8'd7,  9'd261},
{  1'b0, 1'b0,  8'd79,    9'd0},{  1'b0, 1'b0,  8'd78,    9'd0},{  1'b0, 1'b0,  8'd46,  9'd211},{  1'b0, 1'b0,  8'd22,  9'd237},{  1'b0, 1'b1,  8'd10,  9'd326},
{  1'b0, 1'b0,  8'd80,    9'd0},{  1'b0, 1'b0,  8'd79,    9'd0},{  1'b0, 1'b0,  8'd32,  9'd332},{  1'b0, 1'b0,  8'd14,   9'd63},{  1'b0, 1'b1,  8'd10,   9'd97},
{  1'b0, 1'b0,  8'd81,    9'd0},{  1'b0, 1'b0,  8'd80,    9'd0},{  1'b0, 1'b0,  8'd16,  9'd238},{  1'b0, 1'b0,  8'd11,  9'd195},{  1'b0, 1'b1,   8'd5,  9'd339},
{  1'b0, 1'b0,  8'd82,    9'd0},{  1'b0, 1'b0,  8'd81,    9'd0},{  1'b0, 1'b0,  8'd12,  9'd277},{  1'b0, 1'b0,   8'd7,  9'd161},{  1'b0, 1'b1,   8'd1,  9'd185},
{  1'b0, 1'b0,  8'd83,    9'd0},{  1'b0, 1'b0,  8'd82,    9'd0},{  1'b0, 1'b0,  8'd29,  9'd148},{  1'b0, 1'b0,  8'd17,   9'd73},{  1'b0, 1'b1,   8'd3,   9'd66},
{  1'b0, 1'b0,  8'd84,    9'd0},{  1'b0, 1'b0,  8'd83,    9'd0},{  1'b0, 1'b0,  8'd43,  9'd155},{  1'b0, 1'b0,  8'd37,  9'd160},{  1'b0, 1'b1,   8'd9,  9'd192},
{  1'b0, 1'b0,  8'd85,    9'd0},{  1'b0, 1'b0,  8'd84,    9'd0},{  1'b0, 1'b0,  8'd18,  9'd238},{  1'b0, 1'b0,  8'd15,  9'd158},{  1'b0, 1'b1,   8'd6,   9'd37},
{  1'b0, 1'b0,  8'd86,    9'd0},{  1'b0, 1'b0,  8'd85,    9'd0},{  1'b0, 1'b0,   8'd8,  9'd254},{  1'b0, 1'b0,   8'd5,  9'd166},{  1'b0, 1'b1,   8'd0,    9'd4},
{  1'b0, 1'b0,  8'd87,    9'd0},{  1'b0, 1'b0,  8'd86,    9'd0},{  1'b0, 1'b0,  8'd55,   9'd34},{  1'b0, 1'b0,   8'd7,  9'd298},{  1'b0, 1'b1,   8'd2,  9'd107},
{  1'b0, 1'b0,  8'd88,    9'd0},{  1'b0, 1'b0,  8'd87,    9'd0},{  1'b0, 1'b0,  8'd57,  9'd323},{  1'b0, 1'b0,  8'd17,   9'd96},{  1'b0, 1'b1,   8'd4,  9'd213},
{  1'b0, 1'b0,  8'd89,    9'd0},{  1'b0, 1'b0,  8'd88,    9'd0},{  1'b0, 1'b0,  8'd41,  9'd214},{  1'b0, 1'b0,  8'd20,  9'd235},{  1'b0, 1'b1,  8'd13,  9'd187},
{  1'b0, 1'b0,  8'd90,    9'd0},{  1'b0, 1'b0,  8'd89,    9'd0},{  1'b0, 1'b0,  8'd16,  9'd145},{  1'b0, 1'b0,   8'd6,  9'd338},{  1'b0, 1'b1,   8'd1,  9'd274},
{  1'b0, 1'b0,  8'd91,    9'd0},{  1'b0, 1'b0,  8'd90,    9'd0},{  1'b0, 1'b0,  8'd59,  9'd331},{  1'b0, 1'b0,  8'd13,  9'd287},{  1'b0, 1'b1,   8'd4,  9'd299},
{  1'b0, 1'b0,  8'd92,    9'd0},{  1'b0, 1'b0,  8'd91,    9'd0},{  1'b0, 1'b0,  8'd19,  9'd315},{  1'b0, 1'b0,   8'd6,   9'd14},{  1'b0, 1'b1,   8'd5,  9'd242},
{  1'b0, 1'b0,  8'd93,    9'd0},{  1'b0, 1'b0,  8'd92,    9'd0},{  1'b0, 1'b0,  8'd59,  9'd211},{  1'b0, 1'b0,  8'd48,  9'd142},{  1'b0, 1'b1,  8'd33,    9'd5},
{  1'b0, 1'b0,  8'd94,    9'd0},{  1'b0, 1'b0,  8'd93,    9'd0},{  1'b0, 1'b0,  8'd53,  9'd358},{  1'b0, 1'b0,  8'd24,  9'd359},{  1'b0, 1'b1,   8'd3,  9'd296},
{  1'b0, 1'b0,  8'd95,    9'd0},{  1'b0, 1'b0,  8'd94,    9'd0},{  1'b0, 1'b0,  8'd15,   9'd57},{  1'b0, 1'b0,  8'd15,  9'd139},{  1'b0, 1'b1,   8'd5,  9'd300},
{  1'b0, 1'b0,  8'd96,    9'd0},{  1'b0, 1'b0,  8'd95,    9'd0},{  1'b0, 1'b0,  8'd52,  9'd210},{  1'b0, 1'b0,  8'd40,  9'd354},{  1'b0, 1'b1,  8'd18,  9'd126},
{  1'b0, 1'b0,  8'd97,    9'd0},{  1'b0, 1'b0,  8'd96,    9'd0},{  1'b0, 1'b0,  8'd25,  9'd116},{  1'b0, 1'b0,   8'd8,  9'd253},{  1'b0, 1'b1,   8'd8,   9'd28},
{  1'b0, 1'b0,  8'd98,    9'd0},{  1'b0, 1'b0,  8'd97,    9'd0},{  1'b0, 1'b0,   8'd9,  9'd229},{  1'b0, 1'b0,   8'd6,  9'd335},{  1'b0, 1'b1,   8'd0,  9'd154},
{  1'b0, 1'b0,  8'd99,    9'd0},{  1'b0, 1'b0,  8'd98,    9'd0},{  1'b0, 1'b0,  8'd14,  9'd252},{  1'b0, 1'b0,  8'd14,  9'd254},{  1'b0, 1'b1,  8'd11,  9'd202},
{  1'b0, 1'b0, 8'd100,    9'd0},{  1'b0, 1'b0,  8'd99,    9'd0},{  1'b0, 1'b0,  8'd18,   9'd48},{  1'b0, 1'b0,  8'd12,  9'd173},{  1'b0, 1'b1,  8'd10,  9'd126},
{  1'b0, 1'b0, 8'd101,    9'd0},{  1'b0, 1'b0, 8'd100,    9'd0},{  1'b0, 1'b0,  8'd53,   9'd72},{  1'b0, 1'b0,  8'd16,   9'd14},{  1'b0, 1'b1,   8'd2,   9'd85},
{  1'b0, 1'b0, 8'd102,    9'd0},{  1'b0, 1'b0, 8'd101,    9'd0},{  1'b0, 1'b0,  8'd59,   9'd34},{  1'b0, 1'b0,  8'd18,   9'd88},{  1'b0, 1'b1,   8'd7,  9'd102},
{  1'b0, 1'b0, 8'd103,    9'd0},{  1'b0, 1'b0, 8'd102,    9'd0},{  1'b0, 1'b0,  8'd14,  9'd312},{  1'b0, 1'b0,  8'd12,   9'd23},{  1'b0, 1'b1,   8'd4,  9'd100},
{  1'b0, 1'b0, 8'd104,    9'd0},{  1'b0, 1'b0, 8'd103,    9'd0},{  1'b0, 1'b0,  8'd48,   9'd82},{  1'b0, 1'b0,  8'd30,  9'd332},{  1'b0, 1'b1,  8'd18,  9'd181},
{  1'b0, 1'b0, 8'd105,    9'd0},{  1'b0, 1'b0, 8'd104,    9'd0},{  1'b0, 1'b0,  8'd44,  9'd135},{  1'b0, 1'b0,  8'd11,   9'd11},{  1'b0, 1'b1,   8'd5,  9'd136},
{  1'b0, 1'b0, 8'd106,    9'd0},{  1'b0, 1'b0, 8'd105,    9'd0},{  1'b0, 1'b0,  8'd39,   9'd19},{  1'b0, 1'b0,  8'd15,  9'd229},{  1'b0, 1'b1,  8'd10,  9'd112},
{  1'b0, 1'b0, 8'd107,    9'd0},{  1'b0, 1'b0, 8'd106,    9'd0},{  1'b0, 1'b0,  8'd50,  9'd123},{  1'b0, 1'b0,  8'd17,   9'd56},{  1'b0, 1'b1,   8'd0,  9'd174},
{  1'b0, 1'b0, 8'd108,    9'd0},{  1'b0, 1'b0, 8'd107,    9'd0},{  1'b0, 1'b0,  8'd58,   9'd36},{  1'b0, 1'b0,  8'd18,  9'd168},{  1'b0, 1'b1,  8'd12,  9'd344},
{  1'b0, 1'b0, 8'd109,    9'd0},{  1'b0, 1'b0, 8'd108,    9'd0},{  1'b0, 1'b0,  8'd54,  9'd285},{  1'b0, 1'b0,   8'd7,  9'd278},{  1'b0, 1'b1,   8'd2,  9'd145},
{  1'b0, 1'b0, 8'd110,    9'd0},{  1'b0, 1'b0, 8'd109,    9'd0},{  1'b0, 1'b0,  8'd18,  9'd101},{  1'b0, 1'b0,  8'd16,   9'd87},{  1'b0, 1'b1,  8'd12,   9'd66},
{  1'b0, 1'b0, 8'd111,    9'd0},{  1'b0, 1'b0, 8'd110,    9'd0},{  1'b0, 1'b0,  8'd16,  9'd244},{  1'b0, 1'b0,  8'd13,  9'd317},{  1'b0, 1'b1,   8'd0,  9'd213},
{  1'b0, 1'b0, 8'd112,    9'd0},{  1'b0, 1'b0, 8'd111,    9'd0},{  1'b0, 1'b0,  8'd27,   9'd51},{  1'b0, 1'b0,  8'd15,   9'd60},{  1'b0, 1'b1,   8'd2,  9'd286},
{  1'b0, 1'b0, 8'd113,    9'd0},{  1'b0, 1'b0, 8'd112,    9'd0},{  1'b0, 1'b0,  8'd19,  9'd212},{  1'b0, 1'b0,   8'd4,  9'd310},{  1'b0, 1'b1,   8'd0,  9'd267},
{  1'b0, 1'b0, 8'd114,    9'd0},{  1'b0, 1'b0, 8'd113,    9'd0},{  1'b0, 1'b0,  8'd50,  9'd134},{  1'b0, 1'b0,  8'd37,  9'd242},{  1'b0, 1'b1,  8'd29,   9'd84},
{  1'b0, 1'b0, 8'd115,    9'd0},{  1'b0, 1'b0, 8'd114,    9'd0},{  1'b0, 1'b0,  8'd12,   9'd43},{  1'b0, 1'b0,  8'd11,  9'd135},{  1'b0, 1'b1,   8'd8,  9'd281},
{  1'b0, 1'b0, 8'd116,    9'd0},{  1'b0, 1'b0, 8'd115,    9'd0},{  1'b0, 1'b0,  8'd43,  9'd327},{  1'b0, 1'b0,   8'd3,  9'd300},{  1'b0, 1'b1,   8'd1,  9'd315},
{  1'b0, 1'b0, 8'd117,    9'd0},{  1'b0, 1'b0, 8'd116,    9'd0},{  1'b0, 1'b0,  8'd11,  9'd262},{  1'b0, 1'b0,   8'd6,  9'd171},{  1'b0, 1'b1,   8'd3,   9'd45},
{  1'b0, 1'b0, 8'd118,    9'd0},{  1'b0, 1'b0, 8'd117,    9'd0},{  1'b0, 1'b0,  8'd50,  9'd155},{  1'b0, 1'b0,  8'd17,  9'd216},{  1'b0, 1'b1,  8'd10,   9'd31},
{  1'b0, 1'b0, 8'd119,    9'd0},{  1'b0, 1'b0, 8'd118,    9'd0},{  1'b0, 1'b0,  8'd36,   9'd24},{  1'b0, 1'b0,  8'd25,   9'd41},{  1'b0, 1'b1,  8'd20,  9'd207},
{  1'b0, 1'b0, 8'd120,    9'd0},{  1'b0, 1'b0, 8'd119,    9'd0},{  1'b0, 1'b0,  8'd15,  9'd358},{  1'b0, 1'b0,  8'd15,  9'd333},{  1'b0, 1'b1,   8'd8,   9'd42},
{  1'b0, 1'b0, 8'd121,    9'd0},{  1'b0, 1'b0, 8'd120,    9'd0},{  1'b0, 1'b0,  8'd28,  9'd284},{  1'b0, 1'b0,  8'd15,  9'd129},{  1'b0, 1'b1,   8'd7,   9'd77},
{  1'b0, 1'b0, 8'd122,    9'd0},{  1'b0, 1'b0, 8'd121,    9'd0},{  1'b0, 1'b0,  8'd53,  9'd206},{  1'b0, 1'b0,  8'd17,   9'd58},{  1'b0, 1'b1,   8'd2,  9'd213},
{  1'b0, 1'b0, 8'd123,    9'd0},{  1'b0, 1'b0, 8'd122,    9'd0},{  1'b0, 1'b0,  8'd10,  9'd319},{  1'b0, 1'b0,   8'd5,  9'd290},{  1'b0, 1'b1,   8'd4,   9'd59},
{  1'b0, 1'b0, 8'd124,    9'd0},{  1'b0, 1'b0, 8'd123,    9'd0},{  1'b0, 1'b0,  8'd51,  9'd274},{  1'b0, 1'b0,  8'd39,  9'd112},{  1'b0, 1'b1,   8'd2,  9'd138},
{  1'b0, 1'b0, 8'd125,    9'd0},{  1'b0, 1'b0, 8'd124,    9'd0},{  1'b0, 1'b0,  8'd29,  9'd122},{  1'b0, 1'b0,  8'd23,  9'd228},{  1'b0, 1'b1,  8'd10,   9'd35},
{  1'b0, 1'b0, 8'd126,    9'd0},{  1'b0, 1'b0, 8'd125,    9'd0},{  1'b0, 1'b0,  8'd15,  9'd286},{  1'b0, 1'b0,  8'd11,  9'd344},{  1'b0, 1'b1,   8'd5,   9'd92},
{  1'b0, 1'b0, 8'd127,    9'd0},{  1'b0, 1'b0, 8'd126,    9'd0},{  1'b0, 1'b0,  8'd19,  9'd243},{  1'b0, 1'b0,  8'd10,  9'd140},{  1'b0, 1'b1,   8'd4,   9'd98},
{  1'b0, 1'b0, 8'd128,    9'd0},{  1'b0, 1'b0, 8'd127,    9'd0},{  1'b0, 1'b0,  8'd56,  9'd120},{  1'b0, 1'b0,  8'd11,  9'd123},{  1'b0, 1'b1,   8'd8,  9'd201},
{  1'b0, 1'b0, 8'd129,    9'd0},{  1'b0, 1'b0, 8'd128,    9'd0},{  1'b0, 1'b0,  8'd24,  9'd343},{  1'b0, 1'b0,  8'd15,  9'd325},{  1'b0, 1'b1,  8'd10,  9'd218},
{  1'b0, 1'b0, 8'd130,    9'd0},{  1'b0, 1'b0, 8'd129,    9'd0},{  1'b0, 1'b0,  8'd14,  9'd325},{  1'b0, 1'b0,  8'd11,  9'd219},{  1'b0, 1'b1,   8'd4,  9'd340},
{  1'b0, 1'b0, 8'd131,    9'd0},{  1'b0, 1'b0, 8'd130,    9'd0},{  1'b0, 1'b0,  8'd32,  9'd242},{  1'b0, 1'b0,  8'd18,   9'd69},{  1'b0, 1'b1,  8'd17,    9'd3},
{  1'b0, 1'b0, 8'd132,    9'd0},{  1'b0, 1'b0, 8'd131,    9'd0},{  1'b0, 1'b0,  8'd33,  9'd279},{  1'b0, 1'b0,  8'd26,  9'd291},{  1'b0, 1'b1,   8'd4,   9'd82},
{  1'b0, 1'b0, 8'd133,    9'd0},{  1'b0, 1'b0, 8'd132,    9'd0},{  1'b0, 1'b0,  8'd18,  9'd110},{  1'b0, 1'b0,  8'd14,   9'd30},{  1'b0, 1'b1,   8'd3,  9'd115},
{  1'b0, 1'b0, 8'd134,    9'd0},{  1'b0, 1'b0, 8'd133,    9'd0},{  1'b0, 1'b0,  8'd11,   9'd69},{  1'b0, 1'b0,   8'd6,  9'd333},{  1'b0, 1'b1,   8'd1,  9'd121},
{  1'b0, 1'b0, 8'd135,    9'd0},{  1'b0, 1'b0, 8'd134,    9'd0},{  1'b0, 1'b0,  8'd48,  9'd166},{  1'b0, 1'b0,  8'd17,  9'd180},{  1'b0, 1'b1,   8'd3,  9'd243},
{  1'b0, 1'b0, 8'd136,    9'd0},{  1'b0, 1'b0, 8'd135,    9'd0},{  1'b0, 1'b0,  8'd38,  9'd203},{  1'b0, 1'b0,   8'd7,  9'd243},{  1'b0, 1'b1,   8'd5,  9'd329},
{  1'b0, 1'b0, 8'd137,    9'd0},{  1'b0, 1'b0, 8'd136,    9'd0},{  1'b0, 1'b0,  8'd56,  9'd184},{  1'b0, 1'b0,  8'd38,  9'd238},{  1'b0, 1'b1,  8'd37,   9'd44},
{  1'b0, 1'b0, 8'd138,    9'd0},{  1'b0, 1'b0, 8'd137,    9'd0},{  1'b0, 1'b0,  8'd26,   9'd28},{  1'b0, 1'b0,   8'd2,  9'd165},{  1'b0, 1'b1,   8'd1,  9'd184},
{  1'b0, 1'b0, 8'd139,    9'd0},{  1'b0, 1'b0, 8'd138,    9'd0},{  1'b0, 1'b0,  8'd45,  9'd180},{  1'b0, 1'b0,  8'd19,  9'd135},{  1'b0, 1'b1,   8'd0,  9'd311},
{  1'b0, 1'b0, 8'd140,    9'd0},{  1'b0, 1'b0, 8'd139,    9'd0},{  1'b0, 1'b0,  8'd27,  9'd239},{  1'b0, 1'b0,  8'd14,  9'd120},{  1'b0, 1'b1,   8'd4,  9'd144},
{  1'b0, 1'b0, 8'd141,    9'd0},{  1'b0, 1'b0, 8'd140,    9'd0},{  1'b0, 1'b0,  8'd57,  9'd225},{  1'b0, 1'b0,  8'd51,  9'd101},{  1'b0, 1'b1,   8'd1,  9'd258},
{  1'b0, 1'b0, 8'd142,    9'd0},{  1'b0, 1'b0, 8'd141,    9'd0},{  1'b0, 1'b0,  8'd38,   9'd79},{  1'b0, 1'b0,  8'd31,   9'd13},{  1'b0, 1'b1,  8'd24,   9'd50},
{  1'b0, 1'b0, 8'd143,    9'd0},{  1'b0, 1'b0, 8'd142,    9'd0},{  1'b0, 1'b0,  8'd13,   9'd44},{  1'b0, 1'b0,  8'd13,  9'd154},{  1'b0, 1'b1,  8'd11,  9'd238},
{  1'b0, 1'b0, 8'd144,    9'd0},{  1'b0, 1'b0, 8'd143,    9'd0},{  1'b0, 1'b0,  8'd55,  9'd267},{  1'b0, 1'b0,  8'd35,  9'd318},{  1'b0, 1'b1,  8'd18,  9'd286},
{  1'b0, 1'b0, 8'd145,    9'd0},{  1'b0, 1'b0, 8'd144,    9'd0},{  1'b0, 1'b0,  8'd49,  9'd293},{  1'b0, 1'b0,  8'd17,  9'd200},{  1'b0, 1'b1,   8'd6,  9'd159},
{  1'b0, 1'b0, 8'd146,    9'd0},{  1'b0, 1'b0, 8'd145,    9'd0},{  1'b0, 1'b0,  8'd19,   9'd61},{  1'b0, 1'b0,   8'd9,  9'd192},{  1'b0, 1'b1,   8'd9,   9'd24},
{  1'b0, 1'b0, 8'd147,    9'd0},{  1'b0, 1'b0, 8'd146,    9'd0},{  1'b0, 1'b0,  8'd19,  9'd217},{  1'b0, 1'b0,  8'd12,  9'd130},{  1'b0, 1'b1,  8'd12,   9'd53},
{  1'b0, 1'b0, 8'd148,    9'd0},{  1'b0, 1'b0, 8'd147,    9'd0},{  1'b0, 1'b0,  8'd49,  9'd223},{  1'b0, 1'b0,  8'd19,  9'd345},{  1'b0, 1'b1,  8'd19,   9'd58},
{  1'b0, 1'b0, 8'd149,    9'd0},{  1'b0, 1'b0, 8'd148,    9'd0},{  1'b0, 1'b0,   8'd9,  9'd235},{  1'b0, 1'b0,   8'd3,  9'd167},{  1'b0, 1'b1,   8'd2,  9'd103},
{  1'b0, 1'b0, 8'd150,    9'd0},{  1'b0, 1'b0, 8'd149,    9'd0},{  1'b0, 1'b0,  8'd41,  9'd356},{  1'b0, 1'b0,  8'd28,  9'd351},{  1'b0, 1'b1,  8'd14,  9'd166},
{  1'b0, 1'b0, 8'd151,    9'd0},{  1'b0, 1'b0, 8'd150,    9'd0},{  1'b0, 1'b0,  8'd41,  9'd338},{  1'b0, 1'b0,   8'd9,  9'd253},{  1'b0, 1'b1,   8'd7,   9'd26},
{  1'b0, 1'b0, 8'd152,    9'd0},{  1'b0, 1'b0, 8'd151,    9'd0},{  1'b0, 1'b0,  8'd36,   9'd84},{  1'b0, 1'b0,  8'd14,  9'd168},{  1'b0, 1'b1,   8'd0,    9'd8},
{  1'b0, 1'b0, 8'd153,    9'd0},{  1'b0, 1'b0, 8'd152,    9'd0},{  1'b0, 1'b0,  8'd30,  9'd189},{  1'b0, 1'b0,  8'd26,   9'd25},{  1'b0, 1'b1,   8'd1,  9'd127},
{  1'b0, 1'b0, 8'd154,    9'd0},{  1'b0, 1'b0, 8'd153,    9'd0},{  1'b0, 1'b0,  8'd25,  9'd338},{  1'b0, 1'b0,  8'd16,  9'd267},{  1'b0, 1'b1,  8'd10,  9'd127},
{  1'b0, 1'b0, 8'd155,    9'd0},{  1'b0, 1'b0, 8'd154,    9'd0},{  1'b0, 1'b0,  8'd31,  9'd121},{  1'b0, 1'b0,   8'd8,   9'd51},{  1'b0, 1'b1,   8'd5,  9'd295},
{  1'b0, 1'b0, 8'd156,    9'd0},{  1'b0, 1'b0, 8'd155,    9'd0},{  1'b0, 1'b0,  8'd13,  9'd305},{  1'b0, 1'b0,   8'd6,  9'd112},{  1'b0, 1'b1,   8'd4,  9'd182},
{  1'b0, 1'b0, 8'd157,    9'd0},{  1'b0, 1'b0, 8'd156,    9'd0},{  1'b0, 1'b0,  8'd47,    9'd5},{  1'b0, 1'b0,  8'd39,  9'd334},{  1'b0, 1'b1,  8'd13,   9'd10},
{  1'b0, 1'b0, 8'd158,    9'd0},{  1'b0, 1'b0, 8'd157,    9'd0},{  1'b0, 1'b0,  8'd42,  9'd267},{  1'b0, 1'b0,   8'd9,    9'd8},{  1'b0, 1'b1,   8'd6,  9'd117},
{  1'b0, 1'b0, 8'd159,    9'd0},{  1'b0, 1'b0, 8'd158,    9'd0},{  1'b0, 1'b0,  8'd33,   9'd79},{  1'b0, 1'b0,  8'd13,  9'd196},{  1'b0, 1'b1,   8'd8,   9'd80},
{  1'b0, 1'b0, 8'd160,    9'd0},{  1'b0, 1'b0, 8'd159,    9'd0},{  1'b0, 1'b0,   8'd6,  9'd312},{  1'b0, 1'b0,   8'd3,  9'd164},{  1'b0, 1'b1,   8'd3,  9'd124},
{  1'b0, 1'b0, 8'd161,    9'd0},{  1'b0, 1'b0, 8'd160,    9'd0},{  1'b0, 1'b0,  8'd45,   9'd56},{  1'b0, 1'b0,  8'd32,  9'd308},{  1'b0, 1'b1,  8'd28,  9'd341},
{  1'b0, 1'b0, 8'd162,    9'd0},{  1'b0, 1'b0, 8'd161,    9'd0},{  1'b0, 1'b0,  8'd55,  9'd244},{  1'b0, 1'b0,  8'd42,  9'd317},{  1'b0, 1'b1,   8'd6,  9'd130},
{  1'b0, 1'b0, 8'd163,    9'd0},{  1'b0, 1'b0, 8'd162,    9'd0},{  1'b0, 1'b0,  8'd40,  9'd179},{  1'b0, 1'b0,  8'd16,  9'd294},{  1'b0, 1'b1,   8'd0,  9'd290},
{  1'b0, 1'b0, 8'd164,    9'd0},{  1'b0, 1'b0, 8'd163,    9'd0},{  1'b0, 1'b0,  8'd56,   9'd21},{  1'b0, 1'b0,   8'd8,   9'd95},{  1'b0, 1'b1,   8'd1,  9'd155},
{  1'b0, 1'b0, 8'd165,    9'd0},{  1'b0, 1'b0, 8'd164,    9'd0},{  1'b0, 1'b0,   8'd9,   9'd93},{  1'b0, 1'b0,   8'd2,   9'd13},{  1'b0, 1'b1,   8'd1,  9'd124},
{  1'b0, 1'b0, 8'd166,    9'd0},{  1'b0, 1'b0, 8'd165,    9'd0},{  1'b0, 1'b0,  8'd52,  9'd324},{  1'b0, 1'b0,  8'd19,  9'd152},{  1'b0, 1'b1,  8'd12,  9'd115},
{  1'b0, 1'b0, 8'd167,    9'd0},{  1'b0, 1'b0, 8'd166,    9'd0},{  1'b0, 1'b0,  8'd43,  9'd348},{  1'b0, 1'b0,  8'd12,  9'd103},{  1'b0, 1'b1,   8'd9,  9'd123},
{  1'b0, 1'b0, 8'd168,    9'd0},{  1'b0, 1'b0, 8'd167,    9'd0},{  1'b0, 1'b0,  8'd58,  9'd217},{  1'b0, 1'b0,  8'd47,  9'd293},{  1'b0, 1'b1,  8'd20,  9'd332},
{  1'b0, 1'b0, 8'd169,    9'd0},{  1'b0, 1'b0, 8'd168,    9'd0},{  1'b0, 1'b0,  8'd17,  9'd352},{  1'b0, 1'b0,  8'd13,  9'd201},{  1'b0, 1'b1,   8'd3,  9'd166},
{  1'b0, 1'b0, 8'd170,    9'd0},{  1'b0, 1'b0, 8'd169,    9'd0},{  1'b0, 1'b0,  8'd49,   9'd69},{  1'b0, 1'b0,  8'd15,  9'd107},{  1'b0, 1'b1,   8'd7,  9'd238},
{  1'b0, 1'b0, 8'd171,    9'd0},{  1'b0, 1'b0, 8'd170,    9'd0},{  1'b0, 1'b0,  8'd34,  9'd107},{  1'b0, 1'b0,  8'd17,   9'd98},{  1'b0, 1'b1,  8'd14,  9'd331},
{  1'b0, 1'b0, 8'd172,    9'd0},{  1'b0, 1'b0, 8'd171,    9'd0},{  1'b0, 1'b0,  8'd19,  9'd289},{  1'b0, 1'b0,  8'd19,  9'd284},{  1'b0, 1'b1,   8'd4,  9'd242},
{  1'b0, 1'b0, 8'd173,    9'd0},{  1'b0, 1'b0, 8'd172,    9'd0},{  1'b0, 1'b0,  8'd31,  9'd129},{  1'b0, 1'b0,  8'd21,  9'd324},{  1'b0, 1'b1,  8'd16,  9'd332},
{  1'b0, 1'b0, 8'd174,    9'd0},{  1'b0, 1'b0, 8'd173,    9'd0},{  1'b0, 1'b0,  8'd40,   9'd56},{  1'b0, 1'b0,  8'd21,  9'd118},{  1'b0, 1'b1,  8'd13,  9'd347},
{  1'b0, 1'b0, 8'd175,    9'd0},{  1'b0, 1'b0, 8'd174,    9'd0},{  1'b0, 1'b0,  8'd51,   9'd41},{  1'b0, 1'b0,  8'd30,  9'd347},{  1'b0, 1'b1,  8'd12,  9'd197},
{  1'b0, 1'b0, 8'd176,    9'd0},{  1'b0, 1'b0, 8'd175,    9'd0},{  1'b0, 1'b0,   8'd7,   9'd10},{  1'b0, 1'b0,   8'd5,   9'd72},{  1'b0, 1'b1,   8'd1,   9'd96},
{  1'b0, 1'b0, 8'd177,    9'd0},{  1'b0, 1'b0, 8'd176,    9'd0},{  1'b0, 1'b0,  8'd42,  9'd262},{  1'b0, 1'b0,   8'd3,   9'd67},{  1'b0, 1'b1,   8'd3,  9'd176},
{  1'b0, 1'b0, 8'd178,    9'd0},{  1'b0, 1'b0, 8'd177,    9'd0},{  1'b0, 1'b0,   8'd8,  9'd162},{  1'b0, 1'b0,   8'd7,   9'd50},{  1'b0, 1'b1,   8'd1,   9'd56},
{  1'b0, 1'b0, 8'd179,    9'd0},{  1'b0, 1'b0, 8'd178,    9'd0},{  1'b0, 1'b0,  8'd36,  9'd303},{  1'b0, 1'b0,  8'd14,  9'd245},{  1'b0, 1'b1,   8'd2,  9'd296}
};
localparam bit [18 : 0] cLARGE_HS_V_TAB_1BY3_PACKED[cLARGE_HS_TAB_1BY3_PACKED_SIZE] = '{
{8'd179, 1'b0,   10'd0},{8'd179, 1'b1, 10'd595},
{8'd178, 1'b0, 10'd590},{8'd178, 1'b1, 10'd596},
{8'd177, 1'b0, 10'd585},{8'd177, 1'b1, 10'd591},
{8'd176, 1'b0, 10'd580},{8'd176, 1'b1, 10'd586},
{8'd175, 1'b0, 10'd575},{8'd175, 1'b1, 10'd581},
{8'd174, 1'b0, 10'd570},{8'd174, 1'b1, 10'd576},
{8'd173, 1'b0, 10'd565},{8'd173, 1'b1, 10'd571},
{8'd172, 1'b0, 10'd560},{8'd172, 1'b1, 10'd566},
{8'd171, 1'b0, 10'd555},{8'd171, 1'b1, 10'd561},
{8'd170, 1'b0, 10'd550},{8'd170, 1'b1, 10'd556},
{8'd169, 1'b0, 10'd545},{8'd169, 1'b1, 10'd551},
{8'd168, 1'b0, 10'd540},{8'd168, 1'b1, 10'd546},
{8'd167, 1'b0, 10'd535},{8'd167, 1'b1, 10'd541},
{8'd166, 1'b0, 10'd530},{8'd166, 1'b1, 10'd536},
{8'd165, 1'b0, 10'd525},{8'd165, 1'b1, 10'd531},
{8'd164, 1'b0, 10'd520},{8'd164, 1'b1, 10'd526},
{8'd163, 1'b0, 10'd515},{8'd163, 1'b1, 10'd521},
{8'd162, 1'b0, 10'd510},{8'd162, 1'b1, 10'd516},
{8'd161, 1'b0, 10'd505},{8'd161, 1'b1, 10'd511},
{8'd160, 1'b0, 10'd500},{8'd160, 1'b1, 10'd506},
{8'd159, 1'b0, 10'd495},{8'd159, 1'b1, 10'd501},
{8'd158, 1'b0, 10'd490},{8'd158, 1'b1, 10'd496},
{8'd157, 1'b0, 10'd485},{8'd157, 1'b1, 10'd491},
{8'd156, 1'b0, 10'd480},{8'd156, 1'b1, 10'd486},
{8'd155, 1'b0, 10'd475},{8'd155, 1'b1, 10'd481},
{8'd154, 1'b0, 10'd470},{8'd154, 1'b1, 10'd476},
{8'd153, 1'b0, 10'd465},{8'd153, 1'b1, 10'd471},
{8'd152, 1'b0, 10'd460},{8'd152, 1'b1, 10'd466},
{8'd151, 1'b0, 10'd455},{8'd151, 1'b1, 10'd461},
{8'd150, 1'b0, 10'd450},{8'd150, 1'b1, 10'd456},
{8'd149, 1'b0, 10'd445},{8'd149, 1'b1, 10'd451},
{8'd148, 1'b0, 10'd440},{8'd148, 1'b1, 10'd446},
{8'd147, 1'b0, 10'd435},{8'd147, 1'b1, 10'd441},
{8'd146, 1'b0, 10'd430},{8'd146, 1'b1, 10'd436},
{8'd145, 1'b0, 10'd425},{8'd145, 1'b1, 10'd431},
{8'd144, 1'b0, 10'd420},{8'd144, 1'b1, 10'd426},
{8'd143, 1'b0, 10'd415},{8'd143, 1'b1, 10'd421},
{8'd142, 1'b0, 10'd410},{8'd142, 1'b1, 10'd416},
{8'd141, 1'b0, 10'd405},{8'd141, 1'b1, 10'd411},
{8'd140, 1'b0, 10'd400},{8'd140, 1'b1, 10'd406},
{8'd139, 1'b0, 10'd395},{8'd139, 1'b1, 10'd401},
{8'd138, 1'b0, 10'd390},{8'd138, 1'b1, 10'd396},
{8'd137, 1'b0, 10'd385},{8'd137, 1'b1, 10'd391},
{8'd136, 1'b0, 10'd380},{8'd136, 1'b1, 10'd386},
{8'd135, 1'b0, 10'd375},{8'd135, 1'b1, 10'd381},
{8'd134, 1'b0, 10'd370},{8'd134, 1'b1, 10'd376},
{8'd133, 1'b0, 10'd365},{8'd133, 1'b1, 10'd371},
{8'd132, 1'b0, 10'd360},{8'd132, 1'b1, 10'd366},
{8'd131, 1'b0, 10'd355},{8'd131, 1'b1, 10'd361},
{8'd130, 1'b0, 10'd350},{8'd130, 1'b1, 10'd356},
{8'd129, 1'b0, 10'd345},{8'd129, 1'b1, 10'd351},
{8'd128, 1'b0, 10'd340},{8'd128, 1'b1, 10'd346},
{8'd127, 1'b0, 10'd335},{8'd127, 1'b1, 10'd341},
{8'd126, 1'b0, 10'd330},{8'd126, 1'b1, 10'd336},
{8'd125, 1'b0, 10'd325},{8'd125, 1'b1, 10'd331},
{8'd124, 1'b0, 10'd320},{8'd124, 1'b1, 10'd326},
{8'd123, 1'b0, 10'd315},{8'd123, 1'b1, 10'd321},
{8'd122, 1'b0, 10'd310},{8'd122, 1'b1, 10'd316},
{8'd121, 1'b0, 10'd305},{8'd121, 1'b1, 10'd311},
{8'd120, 1'b0, 10'd300},{8'd120, 1'b1, 10'd306},
{8'd119, 1'b0, 10'd295},{8'd119, 1'b1, 10'd301},
{8'd118, 1'b0, 10'd290},{8'd118, 1'b1, 10'd296},
{8'd117, 1'b0, 10'd285},{8'd117, 1'b1, 10'd291},
{8'd116, 1'b0, 10'd280},{8'd116, 1'b1, 10'd286},
{8'd115, 1'b0, 10'd275},{8'd115, 1'b1, 10'd281},
{8'd114, 1'b0, 10'd270},{8'd114, 1'b1, 10'd276},
{8'd113, 1'b0, 10'd265},{8'd113, 1'b1, 10'd271},
{8'd112, 1'b0, 10'd260},{8'd112, 1'b1, 10'd266},
{8'd111, 1'b0, 10'd255},{8'd111, 1'b1, 10'd261},
{8'd110, 1'b0, 10'd250},{8'd110, 1'b1, 10'd256},
{8'd109, 1'b0, 10'd245},{8'd109, 1'b1, 10'd251},
{8'd108, 1'b0, 10'd240},{8'd108, 1'b1, 10'd246},
{8'd107, 1'b0, 10'd235},{8'd107, 1'b1, 10'd241},
{8'd106, 1'b0, 10'd230},{8'd106, 1'b1, 10'd236},
{8'd105, 1'b0, 10'd225},{8'd105, 1'b1, 10'd231},
{8'd104, 1'b0, 10'd220},{8'd104, 1'b1, 10'd226},
{8'd103, 1'b0, 10'd215},{8'd103, 1'b1, 10'd221},
{8'd102, 1'b0, 10'd210},{8'd102, 1'b1, 10'd216},
{8'd101, 1'b0, 10'd205},{8'd101, 1'b1, 10'd211},
{8'd100, 1'b0, 10'd200},{8'd100, 1'b1, 10'd206},
{ 8'd99, 1'b0, 10'd195},{ 8'd99, 1'b1, 10'd201},
{ 8'd98, 1'b0, 10'd190},{ 8'd98, 1'b1, 10'd196},
{ 8'd97, 1'b0, 10'd185},{ 8'd97, 1'b1, 10'd191},
{ 8'd96, 1'b0, 10'd180},{ 8'd96, 1'b1, 10'd186},
{ 8'd95, 1'b0, 10'd175},{ 8'd95, 1'b1, 10'd181},
{ 8'd94, 1'b0, 10'd170},{ 8'd94, 1'b1, 10'd176},
{ 8'd93, 1'b0, 10'd165},{ 8'd93, 1'b1, 10'd171},
{ 8'd92, 1'b0, 10'd160},{ 8'd92, 1'b1, 10'd166},
{ 8'd91, 1'b0, 10'd155},{ 8'd91, 1'b1, 10'd161},
{ 8'd90, 1'b0, 10'd150},{ 8'd90, 1'b1, 10'd156},
{ 8'd89, 1'b0, 10'd145},{ 8'd89, 1'b1, 10'd151},
{ 8'd88, 1'b0, 10'd140},{ 8'd88, 1'b1, 10'd146},
{ 8'd87, 1'b0, 10'd135},{ 8'd87, 1'b1, 10'd141},
{ 8'd86, 1'b0, 10'd130},{ 8'd86, 1'b1, 10'd136},
{ 8'd85, 1'b0, 10'd125},{ 8'd85, 1'b1, 10'd131},
{ 8'd84, 1'b0, 10'd120},{ 8'd84, 1'b1, 10'd126},
{ 8'd83, 1'b0, 10'd115},{ 8'd83, 1'b1, 10'd121},
{ 8'd82, 1'b0, 10'd110},{ 8'd82, 1'b1, 10'd116},
{ 8'd81, 1'b0, 10'd105},{ 8'd81, 1'b1, 10'd111},
{ 8'd80, 1'b0, 10'd100},{ 8'd80, 1'b1, 10'd106},
{ 8'd79, 1'b0,  10'd95},{ 8'd79, 1'b1, 10'd101},
{ 8'd78, 1'b0,  10'd90},{ 8'd78, 1'b1,  10'd96},
{ 8'd77, 1'b0,  10'd85},{ 8'd77, 1'b1,  10'd91},
{ 8'd76, 1'b0,  10'd80},{ 8'd76, 1'b1,  10'd86},
{ 8'd75, 1'b0,  10'd75},{ 8'd75, 1'b1,  10'd81},
{ 8'd74, 1'b0,  10'd70},{ 8'd74, 1'b1,  10'd76},
{ 8'd73, 1'b0,  10'd65},{ 8'd73, 1'b1,  10'd71},
{ 8'd72, 1'b0,  10'd60},{ 8'd72, 1'b1,  10'd66},
{ 8'd71, 1'b0,  10'd55},{ 8'd71, 1'b1,  10'd61},
{ 8'd70, 1'b0,  10'd50},{ 8'd70, 1'b1,  10'd56},
{ 8'd69, 1'b0,  10'd45},{ 8'd69, 1'b1,  10'd51},
{ 8'd68, 1'b0,  10'd40},{ 8'd68, 1'b1,  10'd46},
{ 8'd67, 1'b0,  10'd35},{ 8'd67, 1'b1,  10'd41},
{ 8'd66, 1'b0,  10'd30},{ 8'd66, 1'b1,  10'd36},
{ 8'd65, 1'b0,  10'd25},{ 8'd65, 1'b1,  10'd31},
{ 8'd64, 1'b0,  10'd20},{ 8'd64, 1'b1,  10'd26},
{ 8'd63, 1'b0,  10'd15},{ 8'd63, 1'b1,  10'd21},
{ 8'd62, 1'b0,  10'd10},{ 8'd62, 1'b1,  10'd16},
{ 8'd61, 1'b0,   10'd5},{ 8'd61, 1'b1,  10'd11},
{ 8'd60, 1'b0,   10'd1},{ 8'd60, 1'b1,   10'd6},
{ 8'd59, 1'b0, 10'd157},{ 8'd59, 1'b0, 10'd167},{ 8'd59, 1'b1, 10'd212},
{ 8'd58, 1'b0,  10'd92},{ 8'd58, 1'b0, 10'd242},{ 8'd58, 1'b1, 10'd542},
{ 8'd57, 1'b0,  10'd82},{ 8'd57, 1'b0, 10'd142},{ 8'd57, 1'b1, 10'd407},
{ 8'd56, 1'b0, 10'd342},{ 8'd56, 1'b0, 10'd387},{ 8'd56, 1'b1, 10'd522},
{ 8'd55, 1'b0, 10'd137},{ 8'd55, 1'b0, 10'd422},{ 8'd55, 1'b1, 10'd512},
{ 8'd54, 1'b0,   10'd7},{ 8'd54, 1'b0,  10'd62},{ 8'd54, 1'b1, 10'd247},
{ 8'd53, 1'b0, 10'd172},{ 8'd53, 1'b0, 10'd207},{ 8'd53, 1'b1, 10'd312},
{ 8'd52, 1'b0,  10'd83},{ 8'd52, 1'b0, 10'd182},{ 8'd52, 1'b1, 10'd532},
{ 8'd51, 1'b0, 10'd322},{ 8'd51, 1'b0, 10'd408},{ 8'd51, 1'b1, 10'd577},
{ 8'd50, 1'b0, 10'd237},{ 8'd50, 1'b0, 10'd272},{ 8'd50, 1'b1, 10'd292},
{ 8'd49, 1'b0, 10'd427},{ 8'd49, 1'b0, 10'd442},{ 8'd49, 1'b1, 10'd552},
{ 8'd48, 1'b0, 10'd168},{ 8'd48, 1'b0, 10'd222},{ 8'd48, 1'b1, 10'd377},
{ 8'd47, 1'b0,  10'd37},{ 8'd47, 1'b0, 10'd487},{ 8'd47, 1'b1, 10'd543},
{ 8'd46, 1'b0,   10'd8},{ 8'd46, 1'b0,  10'd17},{ 8'd46, 1'b1,  10'd97},
{ 8'd45, 1'b0,  10'd52},{ 8'd45, 1'b0, 10'd397},{ 8'd45, 1'b1, 10'd507},
{ 8'd44, 1'b0,   10'd2},{ 8'd44, 1'b0,  10'd77},{ 8'd44, 1'b1, 10'd227},
{ 8'd43, 1'b0, 10'd122},{ 8'd43, 1'b0, 10'd282},{ 8'd43, 1'b1, 10'd537},
{ 8'd42, 1'b0, 10'd492},{ 8'd42, 1'b0, 10'd513},{ 8'd42, 1'b1, 10'd587},
{ 8'd41, 1'b0, 10'd147},{ 8'd41, 1'b0, 10'd452},{ 8'd41, 1'b1, 10'd457},
{ 8'd40, 1'b0, 10'd183},{ 8'd40, 1'b0, 10'd517},{ 8'd40, 1'b1, 10'd572},
{ 8'd39, 1'b0, 10'd232},{ 8'd39, 1'b0, 10'd323},{ 8'd39, 1'b1, 10'd488},
{ 8'd38, 1'b0, 10'd382},{ 8'd38, 1'b0, 10'd388},{ 8'd38, 1'b1, 10'd412},
{ 8'd37, 1'b0, 10'd123},{ 8'd37, 1'b0, 10'd273},{ 8'd37, 1'b1, 10'd389},
{ 8'd36, 1'b0, 10'd297},{ 8'd36, 1'b0, 10'd462},{ 8'd36, 1'b1, 10'd597},
{ 8'd35, 1'b0,   10'd9},{ 8'd35, 1'b0,  10'd87},{ 8'd35, 1'b1, 10'd423},
{ 8'd34, 1'b0,  10'd42},{ 8'd34, 1'b0,  10'd88},{ 8'd34, 1'b1, 10'd557},
{ 8'd33, 1'b0, 10'd169},{ 8'd33, 1'b0, 10'd362},{ 8'd33, 1'b1, 10'd497},
{ 8'd32, 1'b0, 10'd102},{ 8'd32, 1'b0, 10'd357},{ 8'd32, 1'b1, 10'd508},
{ 8'd31, 1'b0, 10'd413},{ 8'd31, 1'b0, 10'd477},{ 8'd31, 1'b1, 10'd567},
{ 8'd30, 1'b0, 10'd223},{ 8'd30, 1'b0, 10'd467},{ 8'd30, 1'b1, 10'd578},
{ 8'd29, 1'b0, 10'd117},{ 8'd29, 1'b0, 10'd274},{ 8'd29, 1'b1, 10'd327},
{ 8'd28, 1'b0, 10'd307},{ 8'd28, 1'b0, 10'd453},{ 8'd28, 1'b1, 10'd509},
{ 8'd27, 1'b0,  10'd12},{ 8'd27, 1'b0, 10'd262},{ 8'd27, 1'b1, 10'd402},
{ 8'd26, 1'b0, 10'd363},{ 8'd26, 1'b0, 10'd392},{ 8'd26, 1'b1, 10'd468},
{ 8'd25, 1'b0, 10'd187},{ 8'd25, 1'b0, 10'd298},{ 8'd25, 1'b1, 10'd472},
{ 8'd24, 1'b0, 10'd173},{ 8'd24, 1'b0, 10'd347},{ 8'd24, 1'b1, 10'd414},
{ 8'd23, 1'b0,  10'd22},{ 8'd23, 1'b0,  10'd47},{ 8'd23, 1'b1, 10'd328},
{ 8'd22, 1'b0,  10'd43},{ 8'd22, 1'b0,  10'd72},{ 8'd22, 1'b1,  10'd98},
{ 8'd21, 1'b0,  10'd44},{ 8'd21, 1'b0, 10'd568},{ 8'd21, 1'b1, 10'd573},
{ 8'd20, 1'b0, 10'd148},{ 8'd20, 1'b0, 10'd299},{ 8'd20, 1'b1, 10'd544},
{ 8'd19, 1'b0,  10'd53},{ 8'd19, 1'b0, 10'd162},{ 8'd19, 1'b0, 10'd267},{ 8'd19, 1'b0, 10'd337},{ 8'd19, 1'b0, 10'd398},{ 8'd19, 1'b0, 10'd432},{ 8'd19, 1'b0, 10'd437},{ 8'd19, 1'b0, 10'd443},{ 8'd19, 1'b0, 10'd444},{ 8'd19, 1'b0, 10'd533},{ 8'd19, 1'b0, 10'd562},{ 8'd19, 1'b1, 10'd563},
{ 8'd18, 1'b0,  10'd27},{ 8'd18, 1'b0,  10'd38},{ 8'd18, 1'b0, 10'd127},{ 8'd18, 1'b0, 10'd184},{ 8'd18, 1'b0, 10'd202},{ 8'd18, 1'b0, 10'd213},{ 8'd18, 1'b0, 10'd224},{ 8'd18, 1'b0, 10'd243},{ 8'd18, 1'b0, 10'd252},{ 8'd18, 1'b0, 10'd358},{ 8'd18, 1'b0, 10'd367},{ 8'd18, 1'b1, 10'd424},
{ 8'd17, 1'b0,  10'd28},{ 8'd17, 1'b0,  10'd84},{ 8'd17, 1'b0, 10'd118},{ 8'd17, 1'b0, 10'd143},{ 8'd17, 1'b0, 10'd238},{ 8'd17, 1'b0, 10'd293},{ 8'd17, 1'b0, 10'd313},{ 8'd17, 1'b0, 10'd359},{ 8'd17, 1'b0, 10'd378},{ 8'd17, 1'b0, 10'd428},{ 8'd17, 1'b0, 10'd547},{ 8'd17, 1'b1, 10'd558},
{ 8'd16, 1'b0,  10'd13},{ 8'd16, 1'b0,  10'd48},{ 8'd16, 1'b0,  10'd57},{ 8'd16, 1'b0,  10'd63},{ 8'd16, 1'b0, 10'd107},{ 8'd16, 1'b0, 10'd152},{ 8'd16, 1'b0, 10'd208},{ 8'd16, 1'b0, 10'd253},{ 8'd16, 1'b0, 10'd257},{ 8'd16, 1'b0, 10'd473},{ 8'd16, 1'b0, 10'd518},{ 8'd16, 1'b1, 10'd569},
{ 8'd15, 1'b0,  10'd32},{ 8'd15, 1'b0, 10'd128},{ 8'd15, 1'b0, 10'd177},{ 8'd15, 1'b0, 10'd178},{ 8'd15, 1'b0, 10'd233},{ 8'd15, 1'b0, 10'd263},{ 8'd15, 1'b0, 10'd302},{ 8'd15, 1'b0, 10'd303},{ 8'd15, 1'b0, 10'd308},{ 8'd15, 1'b0, 10'd332},{ 8'd15, 1'b0, 10'd348},{ 8'd15, 1'b1, 10'd553},
{ 8'd14, 1'b0,  10'd64},{ 8'd14, 1'b0, 10'd103},{ 8'd14, 1'b0, 10'd197},{ 8'd14, 1'b0, 10'd198},{ 8'd14, 1'b0, 10'd217},{ 8'd14, 1'b0, 10'd352},{ 8'd14, 1'b0, 10'd368},{ 8'd14, 1'b0, 10'd403},{ 8'd14, 1'b0, 10'd454},{ 8'd14, 1'b0, 10'd463},{ 8'd14, 1'b0, 10'd559},{ 8'd14, 1'b1, 10'd598},
{ 8'd13, 1'b0,  10'd23},{ 8'd13, 1'b0,  10'd89},{ 8'd13, 1'b0, 10'd149},{ 8'd13, 1'b0, 10'd158},{ 8'd13, 1'b0, 10'd258},{ 8'd13, 1'b0, 10'd417},{ 8'd13, 1'b0, 10'd418},{ 8'd13, 1'b0, 10'd482},{ 8'd13, 1'b0, 10'd489},{ 8'd13, 1'b0, 10'd498},{ 8'd13, 1'b0, 10'd548},{ 8'd13, 1'b1, 10'd574},
{ 8'd12, 1'b0,  10'd18},{ 8'd12, 1'b0, 10'd112},{ 8'd12, 1'b0, 10'd203},{ 8'd12, 1'b0, 10'd218},{ 8'd12, 1'b0, 10'd244},{ 8'd12, 1'b0, 10'd254},{ 8'd12, 1'b0, 10'd277},{ 8'd12, 1'b0, 10'd438},{ 8'd12, 1'b0, 10'd439},{ 8'd12, 1'b0, 10'd534},{ 8'd12, 1'b0, 10'd538},{ 8'd12, 1'b1, 10'd579},
{ 8'd11, 1'b0,  10'd67},{ 8'd11, 1'b0,  10'd78},{ 8'd11, 1'b0, 10'd108},{ 8'd11, 1'b0, 10'd199},{ 8'd11, 1'b0, 10'd228},{ 8'd11, 1'b0, 10'd278},{ 8'd11, 1'b0, 10'd287},{ 8'd11, 1'b0, 10'd333},{ 8'd11, 1'b0, 10'd343},{ 8'd11, 1'b0, 10'd353},{ 8'd11, 1'b0, 10'd372},{ 8'd11, 1'b1, 10'd419},
{ 8'd10, 1'b0,  10'd24},{ 8'd10, 1'b0,  10'd68},{ 8'd10, 1'b0,  10'd99},{ 8'd10, 1'b0, 10'd104},{ 8'd10, 1'b0, 10'd204},{ 8'd10, 1'b0, 10'd234},{ 8'd10, 1'b0, 10'd294},{ 8'd10, 1'b0, 10'd317},{ 8'd10, 1'b0, 10'd329},{ 8'd10, 1'b0, 10'd338},{ 8'd10, 1'b0, 10'd349},{ 8'd10, 1'b1, 10'd474},
{  8'd9, 1'b0,  10'd39},{  8'd9, 1'b0,  10'd49},{  8'd9, 1'b0,  10'd58},{  8'd9, 1'b0, 10'd124},{  8'd9, 1'b0, 10'd192},{  8'd9, 1'b0, 10'd433},{  8'd9, 1'b0, 10'd434},{  8'd9, 1'b0, 10'd447},{  8'd9, 1'b0, 10'd458},{  8'd9, 1'b0, 10'd493},{  8'd9, 1'b0, 10'd527},{  8'd9, 1'b1, 10'd539},
{  8'd8, 1'b0,  10'd59},{  8'd8, 1'b0,  10'd93},{  8'd8, 1'b0, 10'd132},{  8'd8, 1'b0, 10'd188},{  8'd8, 1'b0, 10'd189},{  8'd8, 1'b0, 10'd279},{  8'd8, 1'b0, 10'd304},{  8'd8, 1'b0, 10'd344},{  8'd8, 1'b0, 10'd478},{  8'd8, 1'b0, 10'd499},{  8'd8, 1'b0, 10'd523},{  8'd8, 1'b1, 10'd592},
{  8'd7, 1'b0,  10'd79},{  8'd7, 1'b0,  10'd94},{  8'd7, 1'b0, 10'd113},{  8'd7, 1'b0, 10'd138},{  8'd7, 1'b0, 10'd214},{  8'd7, 1'b0, 10'd248},{  8'd7, 1'b0, 10'd309},{  8'd7, 1'b0, 10'd383},{  8'd7, 1'b0, 10'd459},{  8'd7, 1'b0, 10'd554},{  8'd7, 1'b0, 10'd582},{  8'd7, 1'b1, 10'd593},
{  8'd6, 1'b0,  10'd14},{  8'd6, 1'b0, 10'd129},{  8'd6, 1'b0, 10'd153},{  8'd6, 1'b0, 10'd163},{  8'd6, 1'b0, 10'd193},{  8'd6, 1'b0, 10'd288},{  8'd6, 1'b0, 10'd373},{  8'd6, 1'b0, 10'd429},{  8'd6, 1'b0, 10'd483},{  8'd6, 1'b0, 10'd494},{  8'd6, 1'b0, 10'd502},{  8'd6, 1'b1, 10'd514},
{  8'd5, 1'b0,  10'd33},{  8'd5, 1'b0,  10'd34},{  8'd5, 1'b0, 10'd109},{  8'd5, 1'b0, 10'd133},{  8'd5, 1'b0, 10'd164},{  8'd5, 1'b0, 10'd179},{  8'd5, 1'b0, 10'd229},{  8'd5, 1'b0, 10'd318},{  8'd5, 1'b0, 10'd334},{  8'd5, 1'b0, 10'd384},{  8'd5, 1'b0, 10'd479},{  8'd5, 1'b1, 10'd583},
{  8'd4, 1'b0,  10'd29},{  8'd4, 1'b0, 10'd144},{  8'd4, 1'b0, 10'd159},{  8'd4, 1'b0, 10'd219},{  8'd4, 1'b0, 10'd268},{  8'd4, 1'b0, 10'd319},{  8'd4, 1'b0, 10'd339},{  8'd4, 1'b0, 10'd354},{  8'd4, 1'b0, 10'd364},{  8'd4, 1'b0, 10'd404},{  8'd4, 1'b0, 10'd484},{  8'd4, 1'b1, 10'd564},
{  8'd3, 1'b0, 10'd119},{  8'd3, 1'b0, 10'd174},{  8'd3, 1'b0, 10'd283},{  8'd3, 1'b0, 10'd289},{  8'd3, 1'b0, 10'd369},{  8'd3, 1'b0, 10'd379},{  8'd3, 1'b0, 10'd448},{  8'd3, 1'b0, 10'd503},{  8'd3, 1'b0, 10'd504},{  8'd3, 1'b0, 10'd549},{  8'd3, 1'b0, 10'd588},{  8'd3, 1'b1, 10'd589},
{  8'd2, 1'b0,  10'd54},{  8'd2, 1'b0,  10'd73},{  8'd2, 1'b0, 10'd139},{  8'd2, 1'b0, 10'd209},{  8'd2, 1'b0, 10'd249},{  8'd2, 1'b0, 10'd264},{  8'd2, 1'b0, 10'd314},{  8'd2, 1'b0, 10'd324},{  8'd2, 1'b0, 10'd393},{  8'd2, 1'b0, 10'd449},{  8'd2, 1'b0, 10'd528},{  8'd2, 1'b1, 10'd599},
{  8'd1, 1'b0,  10'd19},{  8'd1, 1'b0, 10'd114},{  8'd1, 1'b0, 10'd154},{  8'd1, 1'b0, 10'd284},{  8'd1, 1'b0, 10'd374},{  8'd1, 1'b0, 10'd394},{  8'd1, 1'b0, 10'd409},{  8'd1, 1'b0, 10'd469},{  8'd1, 1'b0, 10'd524},{  8'd1, 1'b0, 10'd529},{  8'd1, 1'b0, 10'd584},{  8'd1, 1'b1, 10'd594},
{  8'd0, 1'b0,   10'd3},{  8'd0, 1'b0,   10'd4},{  8'd0, 1'b0,  10'd69},{  8'd0, 1'b0,  10'd74},{  8'd0, 1'b0, 10'd134},{  8'd0, 1'b0, 10'd194},{  8'd0, 1'b0, 10'd239},{  8'd0, 1'b0, 10'd259},{  8'd0, 1'b0, 10'd269},{  8'd0, 1'b0, 10'd399},{  8'd0, 1'b0, 10'd464},{  8'd0, 1'b1, 10'd519}
};
localparam int          cLARGE_HS_TAB_2BY5_PACKED_SIZE = 648;
localparam bit [18 : 0] cLARGE_HS_TAB_2BY5_PACKED[cLARGE_HS_TAB_2BY5_PACKED_SIZE] = '{
{  1'b1, 1'b0, 8'd179,    9'd1},{  1'b0, 1'b0,  8'd72,    9'd0},{  1'b0, 1'b0,  8'd71,  9'd284},{  1'b0, 1'b0,  8'd32,  9'd263},{  1'b0, 1'b0,   8'd0,   9'd46},{  1'b0, 1'b1,   8'd0,  9'd176},
{  1'b0, 1'b0,  8'd73,    9'd0},{  1'b0, 1'b0,  8'd72,    9'd0},{  1'b0, 1'b0,  8'd45,   9'd66},{  1'b0, 1'b0,  8'd23,  9'd173},{  1'b0, 1'b0,  8'd19,  9'd128},{  1'b0, 1'b1,  8'd17,  9'd243},
{  1'b0, 1'b0,  8'd74,    9'd0},{  1'b0, 1'b0,  8'd73,    9'd0},{  1'b0, 1'b0,  8'd40,  9'd137},{  1'b0, 1'b0,  8'd28,  9'd214},{  1'b0, 1'b0,  8'd11,  9'd355},{  1'b0, 1'b1,   8'd6,  9'd312},
{  1'b0, 1'b0,  8'd75,    9'd0},{  1'b0, 1'b0,  8'd74,    9'd0},{  1'b0, 1'b0,  8'd49,  9'd298},{  1'b0, 1'b0,  8'd23,  9'd213},{  1'b0, 1'b0,  8'd12,  9'd311},{  1'b0, 1'b1,   8'd1,  9'd127},
{  1'b0, 1'b0,  8'd76,    9'd0},{  1'b0, 1'b0,  8'd75,    9'd0},{  1'b0, 1'b0,  8'd71,  9'd137},{  1'b0, 1'b0,  8'd16,  9'd263},{  1'b0, 1'b0,  8'd13,  9'd332},{  1'b0, 1'b1,   8'd5,  9'd189},
{  1'b0, 1'b0,  8'd77,    9'd0},{  1'b0, 1'b0,  8'd76,    9'd0},{  1'b0, 1'b0,  8'd66,  9'd314},{  1'b0, 1'b0,  8'd14,   9'd20},{  1'b0, 1'b0,   8'd5,  9'd103},{  1'b0, 1'b1,   8'd4,  9'd201},
{  1'b0, 1'b0,  8'd78,    9'd0},{  1'b0, 1'b0,  8'd77,    9'd0},{  1'b0, 1'b0,  8'd44,  9'd150},{  1'b0, 1'b0,  8'd17,   9'd54},{  1'b0, 1'b0,  8'd17,  9'd249},{  1'b0, 1'b1,  8'd10,  9'd229},
{  1'b0, 1'b0,  8'd79,    9'd0},{  1'b0, 1'b0,  8'd78,    9'd0},{  1'b0, 1'b0,  8'd61,  9'd317},{  1'b0, 1'b0,  8'd32,   9'd61},{  1'b0, 1'b0,  8'd24,  9'd160},{  1'b0, 1'b1,   8'd9,  9'd312},
{  1'b0, 1'b0,  8'd80,    9'd0},{  1'b0, 1'b0,  8'd79,    9'd0},{  1'b0, 1'b0,  8'd46,   9'd88},{  1'b0, 1'b0,  8'd20,  9'd177},{  1'b0, 1'b0,  8'd12,  9'd135},{  1'b0, 1'b1,   8'd8,  9'd223},
{  1'b0, 1'b0,  8'd81,    9'd0},{  1'b0, 1'b0,  8'd80,    9'd0},{  1'b0, 1'b0,  8'd43,  9'd280},{  1'b0, 1'b0,  8'd19,  9'd219},{  1'b0, 1'b0,  8'd10,    9'd8},{  1'b0, 1'b1,   8'd2,   9'd97},
{  1'b0, 1'b0,  8'd82,    9'd0},{  1'b0, 1'b0,  8'd81,    9'd0},{  1'b0, 1'b0,  8'd67,   9'd99},{  1'b0, 1'b0,  8'd21,  9'd230},{  1'b0, 1'b0,  8'd18,  9'd226},{  1'b0, 1'b1,  8'd11,  9'd144},
{  1'b0, 1'b0,  8'd83,    9'd0},{  1'b0, 1'b0,  8'd82,    9'd0},{  1'b0, 1'b0,  8'd42,  9'd160},{  1'b0, 1'b0,  8'd17,  9'd108},{  1'b0, 1'b0,  8'd15,  9'd166},{  1'b0, 1'b1,  8'd12,   9'd62},
{  1'b0, 1'b0,  8'd84,    9'd0},{  1'b0, 1'b0,  8'd83,    9'd0},{  1'b0, 1'b0,  8'd46,  9'd203},{  1'b0, 1'b0,  8'd21,   9'd38},{  1'b0, 1'b0,   8'd2,  9'd224},{  1'b0, 1'b1,   8'd0,  9'd134},
{  1'b0, 1'b0,  8'd85,    9'd0},{  1'b0, 1'b0,  8'd84,    9'd0},{  1'b0, 1'b0,  8'd60,  9'd205},{  1'b0, 1'b0,   8'd8,  9'd309},{  1'b0, 1'b0,   8'd7,  9'd328},{  1'b0, 1'b1,   8'd0,  9'd137},
{  1'b0, 1'b0,  8'd86,    9'd0},{  1'b0, 1'b0,  8'd85,    9'd0},{  1'b0, 1'b0,  8'd47,  9'd217},{  1'b0, 1'b0,  8'd27,  9'd309},{  1'b0, 1'b0,  8'd26,  9'd289},{  1'b0, 1'b1,  8'd14,  9'd237},
{  1'b0, 1'b0,  8'd87,    9'd0},{  1'b0, 1'b0,  8'd86,    9'd0},{  1'b0, 1'b0,  8'd57,  9'd122},{  1'b0, 1'b0,  8'd23,  9'd354},{  1'b0, 1'b0,  8'd22,  9'd264},{  1'b0, 1'b1,  8'd14,  9'd203},
{  1'b0, 1'b0,  8'd88,    9'd0},{  1'b0, 1'b0,  8'd87,    9'd0},{  1'b0, 1'b0,  8'd59,   9'd97},{  1'b0, 1'b0,  8'd21,  9'd186},{  1'b0, 1'b0,  8'd17,  9'd238},{  1'b0, 1'b1,  8'd15,  9'd245},
{  1'b0, 1'b0,  8'd89,    9'd0},{  1'b0, 1'b0,  8'd88,    9'd0},{  1'b0, 1'b0,  8'd59,   9'd11},{  1'b0, 1'b0,  8'd23,  9'd228},{  1'b0, 1'b0,   8'd8,  9'd324},{  1'b0, 1'b1,   8'd4,  9'd119},
{  1'b0, 1'b0,  8'd90,    9'd0},{  1'b0, 1'b0,  8'd89,    9'd0},{  1'b0, 1'b0,  8'd63,  9'd196},{  1'b0, 1'b0,  8'd21,  9'd112},{  1'b0, 1'b0,   8'd9,  9'd206},{  1'b0, 1'b1,   8'd7,  9'd161},
{  1'b0, 1'b0,  8'd91,    9'd0},{  1'b0, 1'b0,  8'd90,    9'd0},{  1'b0, 1'b0,  8'd68,  9'd122},{  1'b0, 1'b0,  8'd11,  9'd326},{  1'b0, 1'b0,   8'd8,  9'd214},{  1'b0, 1'b1,   8'd6,  9'd335},
{  1'b0, 1'b0,  8'd92,    9'd0},{  1'b0, 1'b0,  8'd91,    9'd0},{  1'b0, 1'b0,  8'd59,   9'd14},{  1'b0, 1'b0,  8'd13,  9'd277},{  1'b0, 1'b0,   8'd5,  9'd166},{  1'b0, 1'b1,   8'd1,  9'd315},
{  1'b0, 1'b0,  8'd93,    9'd0},{  1'b0, 1'b0,  8'd92,    9'd0},{  1'b0, 1'b0,  8'd48,  9'd173},{  1'b0, 1'b0,  8'd22,   9'd13},{  1'b0, 1'b0,  8'd14,  9'd287},{  1'b0, 1'b1,   8'd7,  9'd298},
{  1'b0, 1'b0,  8'd94,    9'd0},{  1'b0, 1'b0,  8'd93,    9'd0},{  1'b0, 1'b0,  8'd56,   9'd70},{  1'b0, 1'b0,  8'd16,   9'd52},{  1'b0, 1'b0,  8'd12,  9'd195},{  1'b0, 1'b1,   8'd2,  9'd107},
{  1'b0, 1'b0,  8'd95,    9'd0},{  1'b0, 1'b0,  8'd94,    9'd0},{  1'b0, 1'b0,  8'd65,  9'd184},{  1'b0, 1'b0,  8'd10,   9'd93},{  1'b0, 1'b0,   8'd9,  9'd254},{  1'b0, 1'b1,   8'd0,    9'd4},
{  1'b0, 1'b0,  8'd96,    9'd0},{  1'b0, 1'b0,  8'd95,    9'd0},{  1'b0, 1'b0,  8'd49,  9'd254},{  1'b0, 1'b0,   8'd5,  9'd242},{  1'b0, 1'b0,   8'd4,   9'd74},{  1'b0, 1'b1,   8'd3,   9'd66},
{  1'b0, 1'b0,  8'd97,    9'd0},{  1'b0, 1'b0,  8'd96,    9'd0},{  1'b0, 1'b0,  8'd56,   9'd98},{  1'b0, 1'b0,  8'd24,  9'd176},{  1'b0, 1'b0,  8'd19,  9'd126},{  1'b0, 1'b1,  8'd16,  9'd158},
{  1'b0, 1'b0,  8'd98,    9'd0},{  1'b0, 1'b0,  8'd97,    9'd0},{  1'b0, 1'b0,  8'd53,  9'd265},{  1'b0, 1'b0,  8'd19,  9'd103},{  1'b0, 1'b0,   8'd8,  9'd141},{  1'b0, 1'b1,   8'd4,  9'd213},
{  1'b0, 1'b0,  8'd99,    9'd0},{  1'b0, 1'b0,  8'd98,    9'd0},{  1'b0, 1'b0,  8'd39,  9'd234},{  1'b0, 1'b0,  8'd22,  9'd285},{  1'b0, 1'b0,  8'd16,   9'd57},{  1'b0, 1'b1,   8'd1,  9'd274},
{  1'b0, 1'b0, 8'd100,    9'd0},{  1'b0, 1'b0,  8'd99,    9'd0},{  1'b0, 1'b0,  8'd50,  9'd279},{  1'b0, 1'b0,  8'd34,   9'd75},{  1'b0, 1'b0,   8'd8,  9'd160},{  1'b0, 1'b1,   8'd6,  9'd333},
{  1'b0, 1'b0, 8'd101,    9'd0},{  1'b0, 1'b0, 8'd100,    9'd0},{  1'b0, 1'b0,  8'd64,  9'd329},{  1'b0, 1'b0,  8'd23,   9'd24},{  1'b0, 1'b0,   8'd4,  9'd299},{  1'b0, 1'b1,   8'd1,  9'd153},
{  1'b0, 1'b0, 8'd102,    9'd0},{  1'b0, 1'b0, 8'd101,    9'd0},{  1'b0, 1'b0,  8'd51,  9'd259},{  1'b0, 1'b0,  8'd18,  9'd329},{  1'b0, 1'b0,   8'd6,  9'd171},{  1'b0, 1'b1,   8'd3,  9'd176},
{  1'b0, 1'b0, 8'd103,    9'd0},{  1'b0, 1'b0, 8'd102,    9'd0},{  1'b0, 1'b0,  8'd53,  9'd182},{  1'b0, 1'b0,  8'd27,  9'd354},{  1'b0, 1'b0,  8'd11,  9'd180},{  1'b0, 1'b1,   8'd6,  9'd143},
{  1'b0, 1'b0, 8'd104,    9'd0},{  1'b0, 1'b0, 8'd103,    9'd0},{  1'b0, 1'b0,  8'd38,  9'd134},{  1'b0, 1'b0,  8'd18,  9'd103},{  1'b0, 1'b0,  8'd15,   9'd63},{  1'b0, 1'b1,   8'd9,   9'd33},
{  1'b0, 1'b0, 8'd105,    9'd0},{  1'b0, 1'b0, 8'd104,    9'd0},{  1'b0, 1'b0,  8'd69,  9'd288},{  1'b0, 1'b0,  8'd31,  9'd209},{  1'b0, 1'b0,  8'd17,  9'd145},{  1'b0, 1'b1,   8'd9,  9'd253},
{  1'b0, 1'b0, 8'd106,    9'd0},{  1'b0, 1'b0, 8'd105,    9'd0},{  1'b0, 1'b0,  8'd57,  9'd248},{  1'b0, 1'b0,  8'd15,  9'd312},{  1'b0, 1'b0,  8'd10,  9'd192},{  1'b0, 1'b1,   8'd0,  9'd154},
{  1'b0, 1'b0, 8'd107,    9'd0},{  1'b0, 1'b0, 8'd106,    9'd0},{  1'b0, 1'b0,  8'd67,  9'd262},{  1'b0, 1'b0,  8'd21,  9'd227},{  1'b0, 1'b0,  8'd13,  9'd100},{  1'b0, 1'b1,   8'd6,  9'd112},
{  1'b0, 1'b0, 8'd108,    9'd0},{  1'b0, 1'b0, 8'd107,    9'd0},{  1'b0, 1'b0,  8'd48,  9'd265},{  1'b0, 1'b0,  8'd17,   9'd87},{  1'b0, 1'b0,  8'd15,  9'd331},{  1'b0, 1'b1,   8'd9,   9'd28},
{  1'b0, 1'b0, 8'd109,    9'd0},{  1'b0, 1'b0, 8'd108,    9'd0},{  1'b0, 1'b0,  8'd65,  9'd107},{  1'b0, 1'b0,  8'd33,  9'd271},{  1'b0, 1'b0,  8'd11,  9'd126},{  1'b0, 1'b1,   8'd2,   9'd85},
{  1'b0, 1'b0, 8'd110,    9'd0},{  1'b0, 1'b0, 8'd109,    9'd0},{  1'b0, 1'b0,  8'd62,  9'd123},{  1'b0, 1'b0,  8'd13,  9'd344},{  1'b0, 1'b0,  8'd12,  9'd202},{  1'b0, 1'b1,   8'd8,  9'd155},
{  1'b0, 1'b0, 8'd111,    9'd0},{  1'b0, 1'b0, 8'd110,    9'd0},{  1'b0, 1'b0,  8'd37,   9'd78},{  1'b0, 1'b0,  8'd13,  9'd173},{  1'b0, 1'b0,  8'd11,  9'd143},{  1'b0, 1'b1,   8'd4,  9'd100},
{  1'b0, 1'b0, 8'd112,    9'd0},{  1'b0, 1'b0, 8'd111,    9'd0},{  1'b0, 1'b0,  8'd50,  9'd293},{  1'b0, 1'b0,  8'd22,  9'd121},{  1'b0, 1'b0,  8'd16,  9'd139},{  1'b0, 1'b1,   8'd7,  9'd102},
{  1'b0, 1'b0, 8'd113,    9'd0},{  1'b0, 1'b0, 8'd112,    9'd0},{  1'b0, 1'b0,  8'd50,  9'd261},{  1'b0, 1'b0,  8'd19,  9'd181},{  1'b0, 1'b0,   8'd5,  9'd136},{  1'b0, 1'b1,   8'd4,  9'd310},
{  1'b0, 1'b0, 8'd114,    9'd0},{  1'b0, 1'b0, 8'd113,    9'd0},{  1'b0, 1'b0,  8'd58,  9'd339},{  1'b0, 1'b0,  8'd18,  9'd105},{  1'b0, 1'b0,  8'd13,  9'd262},{  1'b0, 1'b1,   8'd0,  9'd174},
{  1'b0, 1'b0, 8'd115,    9'd0},{  1'b0, 1'b0, 8'd114,    9'd0},{  1'b0, 1'b0,  8'd68,  9'd202},{  1'b0, 1'b0,  8'd25,  9'd294},{  1'b0, 1'b0,  8'd18,  9'd255},{  1'b0, 1'b1,  8'd11,  9'd112},
{  1'b0, 1'b0, 8'd116,    9'd0},{  1'b0, 1'b0, 8'd115,    9'd0},{  1'b0, 1'b0,  8'd69,   9'd40},{  1'b0, 1'b0,  8'd16,  9'd358},{  1'b0, 1'b0,  8'd15,  9'd161},{  1'b0, 1'b1,   8'd7,  9'd278},
{  1'b0, 1'b0, 8'd117,    9'd0},{  1'b0, 1'b0, 8'd116,    9'd0},{  1'b0, 1'b0,  8'd37,  9'd240},{  1'b0, 1'b0,  8'd13,   9'd23},{  1'b0, 1'b0,  8'd11,   9'd31},{  1'b0, 1'b1,   8'd2,  9'd230},
{  1'b0, 1'b0, 8'd118,    9'd0},{  1'b0, 1'b0, 8'd117,    9'd0},{  1'b0, 1'b0,  8'd58,  9'd147},{  1'b0, 1'b0,  8'd32,    9'd9},{  1'b0, 1'b0,  8'd23,  9'd318},{  1'b0, 1'b1,   8'd0,  9'd213},
{  1'b0, 1'b0, 8'd119,    9'd0},{  1'b0, 1'b0, 8'd118,    9'd0},{  1'b0, 1'b0,  8'd68,  9'd195},{  1'b0, 1'b0,  8'd19,   9'd48},{  1'b0, 1'b0,  8'd14,  9'd317},{  1'b0, 1'b1,   8'd6,   9'd65},
{  1'b0, 1'b0, 8'd120,    9'd0},{  1'b0, 1'b0, 8'd119,    9'd0},{  1'b0, 1'b0,  8'd41,   9'd72},{  1'b0, 1'b0,  8'd21,  9'd345},{  1'b0, 1'b0,   8'd2,  9'd286},{  1'b0, 1'b1,   8'd0,  9'd267},
{  1'b0, 1'b0, 8'd121,    9'd0},{  1'b0, 1'b0, 8'd120,    9'd0},{  1'b0, 1'b0,  8'd37,  9'd123},{  1'b0, 1'b0,  8'd20,  9'd315},{  1'b0, 1'b0,  8'd11,  9'd319},{  1'b0, 1'b1,   8'd3,   9'd67},
{  1'b0, 1'b0, 8'd122,    9'd0},{  1'b0, 1'b0, 8'd121,    9'd0},{  1'b0, 1'b0,  8'd52,  9'd123},{  1'b0, 1'b0,  8'd23,   9'd84},{  1'b0, 1'b0,   8'd3,  9'd167},{  1'b0, 1'b1,   8'd1,  9'd124},
{  1'b0, 1'b0, 8'd123,    9'd0},{  1'b0, 1'b0, 8'd122,    9'd0},{  1'b0, 1'b0,  8'd44,   9'd19},{  1'b0, 1'b0,  8'd34,  9'd187},{  1'b0, 1'b0,  8'd13,   9'd43},{  1'b0, 1'b1,   8'd3,  9'd201},
{  1'b0, 1'b0, 8'd124,    9'd0},{  1'b0, 1'b0, 8'd123,    9'd0},{  1'b0, 1'b0,  8'd69,   9'd44},{  1'b0, 1'b0,  8'd27,  9'd230},{  1'b0, 1'b0,  8'd12,  9'd344},{  1'b0, 1'b1,   8'd9,  9'd281},
{  1'b0, 1'b0, 8'd125,    9'd0},{  1'b0, 1'b0, 8'd124,    9'd0},{  1'b0, 1'b0,  8'd62,  9'd327},{  1'b0, 1'b0,  8'd22,  9'd129},{  1'b0, 1'b0,  8'd18,   9'd65},{  1'b0, 1'b1,  8'd17,  9'd244},
{  1'b0, 1'b0, 8'd126,    9'd0},{  1'b0, 1'b0, 8'd125,    9'd0},{  1'b0, 1'b0,  8'd38,  9'd182},{  1'b0, 1'b0,  8'd13,   9'd66},{  1'b0, 1'b0,   8'd9,   9'd42},{  1'b0, 1'b1,   8'd6,   9'd14},
{  1'b0, 1'b0, 8'd127,    9'd0},{  1'b0, 1'b0, 8'd126,    9'd0},{  1'b0, 1'b0,  8'd57,   9'd96},{  1'b0, 1'b0,  8'd19,  9'd168},{  1'b0, 1'b0,  8'd18,  9'd350},{  1'b0, 1'b1,   8'd8,  9'd208},
{  1'b0, 1'b0, 8'd128,    9'd0},{  1'b0, 1'b0, 8'd127,    9'd0},{  1'b0, 1'b0,  8'd52,  9'd116},{  1'b0, 1'b0,  8'd25,  9'd112},{  1'b0, 1'b0,   8'd8,   9'd48},{  1'b0, 1'b1,   8'd7,   9'd77},
{  1'b0, 1'b0, 8'd129,    9'd0},{  1'b0, 1'b0, 8'd128,    9'd0},{  1'b0, 1'b0,  8'd64,  9'd161},{  1'b0, 1'b0,  8'd22,  9'd332},{  1'b0, 1'b0,  8'd16,  9'd325},{  1'b0, 1'b1,  8'd12,  9'd219},
{  1'b0, 1'b0, 8'd130,    9'd0},{  1'b0, 1'b0, 8'd129,    9'd0},{  1'b0, 1'b0,  8'd47,  9'd312},{  1'b0, 1'b0,  8'd10,  9'd290},{  1'b0, 1'b0,   8'd2,  9'd138},{  1'b0, 1'b1,   8'd2,  9'd213},
{  1'b0, 1'b0, 8'd131,    9'd0},{  1'b0, 1'b0, 8'd130,    9'd0},{  1'b0, 1'b0,  8'd51,   9'd78},{  1'b0, 1'b0,  8'd35,  9'd247},{  1'b0, 1'b0,  8'd12,   9'd69},{  1'b0, 1'b1,   8'd9,  9'd201},
{  1'b0, 1'b0, 8'd132,    9'd0},{  1'b0, 1'b0, 8'd131,    9'd0},{  1'b0, 1'b0,  8'd41,   9'd11},{  1'b0, 1'b0,  8'd33,  9'd184},{  1'b0, 1'b0,  8'd11,   9'd35},{  1'b0, 1'b1,   8'd5,  9'd290},
{  1'b0, 1'b0, 8'd133,    9'd0},{  1'b0, 1'b0, 8'd132,    9'd0},{  1'b0, 1'b0,  8'd46,  9'd359},{  1'b0, 1'b0,  8'd20,  9'd212},{  1'b0, 1'b0,  8'd14,  9'd285},{  1'b0, 1'b1,  8'd11,  9'd140},
{  1'b0, 1'b0, 8'd134,    9'd0},{  1'b0, 1'b0, 8'd133,    9'd0},{  1'b0, 1'b0,  8'd40,  9'd236},{  1'b0, 1'b0,  8'd23,  9'd199},{  1'b0, 1'b0,   8'd6,   9'd37},{  1'b0, 1'b1,   8'd4,   9'd98},
{  1'b0, 1'b0, 8'd135,    9'd0},{  1'b0, 1'b0, 8'd134,    9'd0},{  1'b0, 1'b0,  8'd66,  9'd311},{  1'b0, 1'b0,  8'd22,  9'd353},{  1'b0, 1'b0,  8'd19,  9'd110},{  1'b0, 1'b1,  8'd18,  9'd319},
{  1'b0, 1'b0, 8'd136,    9'd0},{  1'b0, 1'b0, 8'd135,    9'd0},{  1'b0, 1'b0,  8'd45,  9'd181},{  1'b0, 1'b0,  8'd19,   9'd69},{  1'b0, 1'b0,   8'd5,   9'd92},{  1'b0, 1'b1,   8'd4,  9'd340},
{  1'b0, 1'b0, 8'd137,    9'd0},{  1'b0, 1'b0, 8'd136,    9'd0},{  1'b0, 1'b0,  8'd51,  9'd141},{  1'b0, 1'b0,  8'd29,  9'd335},{  1'b0, 1'b0,  8'd16,  9'd333},{  1'b0, 1'b1,   8'd5,  9'd329},
{  1'b0, 1'b0, 8'd138,    9'd0},{  1'b0, 1'b0, 8'd137,    9'd0},{  1'b0, 1'b0,  8'd58,  9'd198},{  1'b0, 1'b0,  8'd16,  9'd129},{  1'b0, 1'b0,  8'd12,  9'd123},{  1'b0, 1'b1,   8'd3,  9'd115},
{  1'b0, 1'b0, 8'd139,    9'd0},{  1'b0, 1'b0, 8'd138,    9'd0},{  1'b0, 1'b0,  8'd36,  9'd275},{  1'b0, 1'b0,  8'd30,    9'd1},{  1'b0, 1'b0,   8'd8,  9'd190},{  1'b0, 1'b1,   8'd1,  9'd184},
{  1'b0, 1'b0, 8'd140,    9'd0},{  1'b0, 1'b0, 8'd139,    9'd0},{  1'b0, 1'b0,  8'd42,  9'd285},{  1'b0, 1'b0,  8'd33,   9'd32},{  1'b0, 1'b0,  8'd16,  9'd337},{  1'b0, 1'b1,   8'd4,  9'd144},
{  1'b0, 1'b0, 8'd141,    9'd0},{  1'b0, 1'b0, 8'd140,    9'd0},{  1'b0, 1'b0,  8'd49,  9'd210},{  1'b0, 1'b0,  8'd35,  9'd336},{  1'b0, 1'b0,  8'd19,  9'd101},{  1'b0, 1'b1,   8'd7,  9'd243},
{  1'b0, 1'b0, 8'd142,    9'd0},{  1'b0, 1'b0, 8'd141,    9'd0},{  1'b0, 1'b0,  8'd42,   9'd49},{  1'b0, 1'b0,  8'd19,  9'd329},{  1'b0, 1'b0,   8'd8,    9'd6},{  1'b0, 1'b1,   8'd1,  9'd123},
{  1'b0, 1'b0, 8'd143,    9'd0},{  1'b0, 1'b0, 8'd142,    9'd0},{  1'b0, 1'b0,  8'd54,   9'd41},{  1'b0, 1'b0,  8'd23,   9'd54},{  1'b0, 1'b0,  8'd11,  9'd218},{  1'b0, 1'b1,   8'd0,  9'd311},
{  1'b0, 1'b0, 8'd144,    9'd0},{  1'b0, 1'b0, 8'd143,    9'd0},{  1'b0, 1'b0,  8'd55,  9'd110},{  1'b0, 1'b0,  8'd21,  9'd237},{  1'b0, 1'b0,  8'd18,  9'd164},{  1'b0, 1'b1,   8'd2,  9'd165},
{  1'b0, 1'b0, 8'd145,    9'd0},{  1'b0, 1'b0, 8'd144,    9'd0},{  1'b0, 1'b0,  8'd43,  9'd250},{  1'b0, 1'b0,  8'd20,  9'd243},{  1'b0, 1'b0,   8'd8,   9'd49},{  1'b0, 1'b1,   8'd1,  9'd155},
{  1'b0, 1'b0, 8'd146,    9'd0},{  1'b0, 1'b0, 8'd145,    9'd0},{  1'b0, 1'b0,  8'd53,   9'd23},{  1'b0, 1'b0,  8'd31,  9'd135},{  1'b0, 1'b0,  8'd12,  9'd238},{  1'b0, 1'b1,  8'd12,   9'd92},
{  1'b0, 1'b0, 8'd147,    9'd0},{  1'b0, 1'b0, 8'd146,    9'd0},{  1'b0, 1'b0,  8'd48,  9'd167},{  1'b0, 1'b0,  8'd30,   9'd66},{  1'b0, 1'b0,  8'd29,   9'd97},{  1'b0, 1'b1,  8'd18,   9'd73},
{  1'b0, 1'b0, 8'd148,    9'd0},{  1'b0, 1'b0, 8'd147,    9'd0},{  1'b0, 1'b0,  8'd38,  9'd340},{  1'b0, 1'b0,  8'd24,  9'd252},{  1'b0, 1'b0,  8'd15,  9'd252},{  1'b0, 1'b1,   8'd3,  9'd229},
{  1'b0, 1'b0, 8'd149,    9'd0},{  1'b0, 1'b0, 8'd148,    9'd0},{  1'b0, 1'b0,  8'd70,   9'd51},{  1'b0, 1'b0,  8'd31,  9'd353},{  1'b0, 1'b0,  8'd22,  9'd300},{  1'b0, 1'b1,  8'd21,  9'd133},
{  1'b0, 1'b0, 8'd150,    9'd0},{  1'b0, 1'b0, 8'd149,    9'd0},{  1'b0, 1'b0,  8'd70,   9'd44},{  1'b0, 1'b0,  8'd14,  9'd154},{  1'b0, 1'b0,  8'd13,   9'd53},{  1'b0, 1'b1,  8'd10,   9'd63},
{  1'b0, 1'b0, 8'd151,    9'd0},{  1'b0, 1'b0, 8'd150,    9'd0},{  1'b0, 1'b0,  8'd71,  9'd156},{  1'b0, 1'b0,  8'd18,  9'd349},{  1'b0, 1'b0,  8'd12,  9'd262},{  1'b0, 1'b1,   8'd3,  9'd166},
{  1'b0, 1'b0, 8'd152,    9'd0},{  1'b0, 1'b0, 8'd151,    9'd0},{  1'b0, 1'b0,  8'd61,   9'd47},{  1'b0, 1'b0,   8'd7,   9'd26},{  1'b0, 1'b0,   8'd7,  9'd344},{  1'b0, 1'b1,   8'd2,  9'd103},
{  1'b0, 1'b0, 8'd153,    9'd0},{  1'b0, 1'b0, 8'd152,    9'd0},{  1'b0, 1'b0,  8'd63,   9'd13},{  1'b0, 1'b0,  8'd22,   9'd79},{  1'b0, 1'b0,  8'd19,  9'd286},{  1'b0, 1'b1,  8'd10,   9'd24},
{  1'b0, 1'b0, 8'd154,    9'd0},{  1'b0, 1'b0, 8'd153,    9'd0},{  1'b0, 1'b0,  8'd39,   9'd67},{  1'b0, 1'b0,  8'd23,  9'd303},{  1'b0, 1'b0,  8'd20,   9'd61},{  1'b0, 1'b1,  8'd20,  9'd217},
{  1'b0, 1'b0, 8'd155,    9'd0},{  1'b0, 1'b0, 8'd154,    9'd0},{  1'b0, 1'b0,  8'd67,  9'd185},{  1'b0, 1'b0,  8'd10,  9'd235},{  1'b0, 1'b0,   8'd5,  9'd295},{  1'b0, 1'b1,   8'd0,    9'd8},
{  1'b0, 1'b0, 8'd156,    9'd0},{  1'b0, 1'b0, 8'd155,    9'd0},{  1'b0, 1'b0,  8'd52,  9'd137},{  1'b0, 1'b0,  8'd20,  9'd345},{  1'b0, 1'b0,  8'd20,   9'd58},{  1'b0, 1'b1,   8'd1,   9'd56},
{  1'b0, 1'b0, 8'd157,    9'd0},{  1'b0, 1'b0, 8'd156,    9'd0},{  1'b0, 1'b0,  8'd65,  9'd306},{  1'b0, 1'b0,  8'd18,  9'd200},{  1'b0, 1'b0,  8'd10,  9'd253},{  1'b0, 1'b1,   8'd6,  9'd130},
{  1'b0, 1'b0, 8'd158,    9'd0},{  1'b0, 1'b0, 8'd157,    9'd0},{  1'b0, 1'b0,  8'd60,  9'd337},{  1'b0, 1'b0,  8'd15,  9'd151},{  1'b0, 1'b0,  8'd14,  9'd305},{  1'b0, 1'b1,  8'd10,   9'd64},
{  1'b0, 1'b0, 8'd159,    9'd0},{  1'b0, 1'b0, 8'd158,    9'd0},{  1'b0, 1'b0,  8'd66,   9'd72},{  1'b0, 1'b0,  8'd28,  9'd351},{  1'b0, 1'b0,  8'd20,  9'd186},{  1'b0, 1'b1,  8'd17,  9'd267},
{  1'b0, 1'b0, 8'd160,    9'd0},{  1'b0, 1'b0, 8'd159,    9'd0},{  1'b0, 1'b0,  8'd36,  9'd125},{  1'b0, 1'b0,  8'd26,  9'd112},{  1'b0, 1'b0,   8'd9,   9'd51},{  1'b0, 1'b1,   8'd4,  9'd182},
{  1'b0, 1'b0, 8'd161,    9'd0},{  1'b0, 1'b0, 8'd160,    9'd0},{  1'b0, 1'b0,  8'd55,   9'd77},{  1'b0, 1'b0,  8'd23,  9'd252},{  1'b0, 1'b0,  8'd10,  9'd101},{  1'b0, 1'b1,   8'd6,  9'd117},
{  1'b0, 1'b0, 8'd162,    9'd0},{  1'b0, 1'b0, 8'd161,    9'd0},{  1'b0, 1'b0,  8'd55,  9'd262},{  1'b0, 1'b0,  8'd15,  9'd213},{  1'b0, 1'b0,   8'd6,  9'd338},{  1'b0, 1'b1,   8'd3,  9'd300},
{  1'b0, 1'b0, 8'd163,    9'd0},{  1'b0, 1'b0, 8'd162,    9'd0},{  1'b0, 1'b0,  8'd36,   9'd69},{  1'b0, 1'b0,  8'd30,  9'd327},{  1'b0, 1'b0,  8'd14,  9'd196},{  1'b0, 1'b1,   8'd3,  9'd124},
{  1'b0, 1'b0, 8'd164,    9'd0},{  1'b0, 1'b0, 8'd163,    9'd0},{  1'b0, 1'b0,  8'd54,  9'd243},{  1'b0, 1'b0,  8'd25,  9'd238},{  1'b0, 1'b0,   8'd9,   9'd80},{  1'b0, 1'b1,   8'd5,  9'd308},
{  1'b0, 1'b0, 8'd165,    9'd0},{  1'b0, 1'b0, 8'd164,    9'd0},{  1'b0, 1'b0,  8'd70,   9'd18},{  1'b0, 1'b0,  8'd22,  9'd198},{  1'b0, 1'b0,  8'd16,  9'd153},{  1'b0, 1'b1,   8'd0,  9'd290},
{  1'b0, 1'b0, 8'd166,    9'd0},{  1'b0, 1'b0, 8'd165,    9'd0},{  1'b0, 1'b0,  8'd45,  9'd296},{  1'b0, 1'b0,  8'd20,  9'd152},{  1'b0, 1'b0,  8'd13,  9'd115},{  1'b0, 1'b1,   8'd1,  9'd258},
{  1'b0, 1'b0, 8'd167,    9'd0},{  1'b0, 1'b0, 8'd166,    9'd0},{  1'b0, 1'b0,  8'd60,  9'd282},{  1'b0, 1'b0,  8'd14,   9'd10},{  1'b0, 1'b0,  8'd10,  9'd123},{  1'b0, 1'b1,   8'd2,   9'd13},
{  1'b0, 1'b0, 8'd168,    9'd0},{  1'b0, 1'b0, 8'd167,    9'd0},{  1'b0, 1'b0,  8'd43,  9'd267},{  1'b0, 1'b0,  8'd28,  9'd275},{  1'b0, 1'b0,  8'd26,  9'd324},{  1'b0, 1'b1,  8'd23,  9'd245},
{  1'b0, 1'b0, 8'd169,    9'd0},{  1'b0, 1'b0, 8'd168,    9'd0},{  1'b0, 1'b0,  8'd56,    9'd8},{  1'b0, 1'b0,  8'd21,  9'd194},{  1'b0, 1'b0,  8'd20,   9'd81},{  1'b0, 1'b1,   8'd3,   9'd45},
{  1'b0, 1'b0, 8'd170,    9'd0},{  1'b0, 1'b0, 8'd169,    9'd0},{  1'b0, 1'b0,  8'd61,  9'd104},{  1'b0, 1'b0,  8'd35,  9'd166},{  1'b0, 1'b0,  8'd17,   9'd74},{  1'b0, 1'b1,   8'd7,  9'd238},
{  1'b0, 1'b0, 8'd171,    9'd0},{  1'b0, 1'b0, 8'd170,    9'd0},{  1'b0, 1'b0,  8'd40,  9'd324},{  1'b0, 1'b0,  8'd17,  9'd294},{  1'b0, 1'b0,  8'd16,  9'd107},{  1'b0, 1'b1,  8'd14,  9'd201},
{  1'b0, 1'b0, 8'd172,    9'd0},{  1'b0, 1'b0, 8'd171,    9'd0},{  1'b0, 1'b0,  8'd39,   9'd41},{  1'b0, 1'b0,  8'd29,  9'd317},{  1'b0, 1'b0,  8'd15,  9'd177},{  1'b0, 1'b1,   8'd4,  9'd242},
{  1'b0, 1'b0, 8'd173,    9'd0},{  1'b0, 1'b0, 8'd172,    9'd0},{  1'b0, 1'b0,  8'd47,  9'd331},{  1'b0, 1'b0,  8'd21,  9'd323},{  1'b0, 1'b0,  8'd17,  9'd342},{  1'b0, 1'b1,  8'd15,  9'd168},
{  1'b0, 1'b0, 8'd174,    9'd0},{  1'b0, 1'b0, 8'd173,    9'd0},{  1'b0, 1'b0,  8'd44,  9'd120},{  1'b0, 1'b0,  8'd20,  9'd284},{  1'b0, 1'b0,  8'd14,  9'd347},{  1'b0, 1'b1,   8'd5,  9'd257},
{  1'b0, 1'b0, 8'd175,    9'd0},{  1'b0, 1'b0, 8'd174,    9'd0},{  1'b0, 1'b0,  8'd54,   9'd57},{  1'b0, 1'b0,  8'd21,   9'd27},{  1'b0, 1'b0,  8'd21,  9'd228},{  1'b0, 1'b1,  8'd13,  9'd197},
{  1'b0, 1'b0, 8'd176,    9'd0},{  1'b0, 1'b0, 8'd175,    9'd0},{  1'b0, 1'b0,  8'd62,  9'd264},{  1'b0, 1'b0,  8'd22,  9'd308},{  1'b0, 1'b0,   8'd7,   9'd10},{  1'b0, 1'b1,   8'd1,  9'd121},
{  1'b0, 1'b0, 8'd177,    9'd0},{  1'b0, 1'b0, 8'd176,    9'd0},{  1'b0, 1'b0,  8'd64,  9'd217},{  1'b0, 1'b0,  8'd34,  9'd293},{  1'b0, 1'b0,  8'd22,  9'd242},{  1'b0, 1'b1,   8'd3,  9'd296},
{  1'b0, 1'b0, 8'd178,    9'd0},{  1'b0, 1'b0, 8'd177,    9'd0},{  1'b0, 1'b0,  8'd63,   9'd82},{  1'b0, 1'b0,   8'd9,  9'd162},{  1'b0, 1'b0,   8'd5,   9'd72},{  1'b0, 1'b1,   8'd1,  9'd185},
{  1'b0, 1'b0, 8'd179,    9'd0},{  1'b0, 1'b0, 8'd178,    9'd0},{  1'b0, 1'b0,  8'd41,    9'd1},{  1'b0, 1'b0,  8'd15,  9'd254},{  1'b0, 1'b0,   8'd7,   9'd50},{  1'b0, 1'b1,   8'd2,  9'd296}
};
localparam bit [18 : 0] cLARGE_HS_V_TAB_2BY5_PACKED[cLARGE_HS_TAB_2BY5_PACKED_SIZE] = '{
{8'd179, 1'b0,   10'd0},{8'd179, 1'b1, 10'd642},
{8'd178, 1'b0, 10'd636},{8'd178, 1'b1, 10'd643},
{8'd177, 1'b0, 10'd630},{8'd177, 1'b1, 10'd637},
{8'd176, 1'b0, 10'd624},{8'd176, 1'b1, 10'd631},
{8'd175, 1'b0, 10'd618},{8'd175, 1'b1, 10'd625},
{8'd174, 1'b0, 10'd612},{8'd174, 1'b1, 10'd619},
{8'd173, 1'b0, 10'd606},{8'd173, 1'b1, 10'd613},
{8'd172, 1'b0, 10'd600},{8'd172, 1'b1, 10'd607},
{8'd171, 1'b0, 10'd594},{8'd171, 1'b1, 10'd601},
{8'd170, 1'b0, 10'd588},{8'd170, 1'b1, 10'd595},
{8'd169, 1'b0, 10'd582},{8'd169, 1'b1, 10'd589},
{8'd168, 1'b0, 10'd576},{8'd168, 1'b1, 10'd583},
{8'd167, 1'b0, 10'd570},{8'd167, 1'b1, 10'd577},
{8'd166, 1'b0, 10'd564},{8'd166, 1'b1, 10'd571},
{8'd165, 1'b0, 10'd558},{8'd165, 1'b1, 10'd565},
{8'd164, 1'b0, 10'd552},{8'd164, 1'b1, 10'd559},
{8'd163, 1'b0, 10'd546},{8'd163, 1'b1, 10'd553},
{8'd162, 1'b0, 10'd540},{8'd162, 1'b1, 10'd547},
{8'd161, 1'b0, 10'd534},{8'd161, 1'b1, 10'd541},
{8'd160, 1'b0, 10'd528},{8'd160, 1'b1, 10'd535},
{8'd159, 1'b0, 10'd522},{8'd159, 1'b1, 10'd529},
{8'd158, 1'b0, 10'd516},{8'd158, 1'b1, 10'd523},
{8'd157, 1'b0, 10'd510},{8'd157, 1'b1, 10'd517},
{8'd156, 1'b0, 10'd504},{8'd156, 1'b1, 10'd511},
{8'd155, 1'b0, 10'd498},{8'd155, 1'b1, 10'd505},
{8'd154, 1'b0, 10'd492},{8'd154, 1'b1, 10'd499},
{8'd153, 1'b0, 10'd486},{8'd153, 1'b1, 10'd493},
{8'd152, 1'b0, 10'd480},{8'd152, 1'b1, 10'd487},
{8'd151, 1'b0, 10'd474},{8'd151, 1'b1, 10'd481},
{8'd150, 1'b0, 10'd468},{8'd150, 1'b1, 10'd475},
{8'd149, 1'b0, 10'd462},{8'd149, 1'b1, 10'd469},
{8'd148, 1'b0, 10'd456},{8'd148, 1'b1, 10'd463},
{8'd147, 1'b0, 10'd450},{8'd147, 1'b1, 10'd457},
{8'd146, 1'b0, 10'd444},{8'd146, 1'b1, 10'd451},
{8'd145, 1'b0, 10'd438},{8'd145, 1'b1, 10'd445},
{8'd144, 1'b0, 10'd432},{8'd144, 1'b1, 10'd439},
{8'd143, 1'b0, 10'd426},{8'd143, 1'b1, 10'd433},
{8'd142, 1'b0, 10'd420},{8'd142, 1'b1, 10'd427},
{8'd141, 1'b0, 10'd414},{8'd141, 1'b1, 10'd421},
{8'd140, 1'b0, 10'd408},{8'd140, 1'b1, 10'd415},
{8'd139, 1'b0, 10'd402},{8'd139, 1'b1, 10'd409},
{8'd138, 1'b0, 10'd396},{8'd138, 1'b1, 10'd403},
{8'd137, 1'b0, 10'd390},{8'd137, 1'b1, 10'd397},
{8'd136, 1'b0, 10'd384},{8'd136, 1'b1, 10'd391},
{8'd135, 1'b0, 10'd378},{8'd135, 1'b1, 10'd385},
{8'd134, 1'b0, 10'd372},{8'd134, 1'b1, 10'd379},
{8'd133, 1'b0, 10'd366},{8'd133, 1'b1, 10'd373},
{8'd132, 1'b0, 10'd360},{8'd132, 1'b1, 10'd367},
{8'd131, 1'b0, 10'd354},{8'd131, 1'b1, 10'd361},
{8'd130, 1'b0, 10'd348},{8'd130, 1'b1, 10'd355},
{8'd129, 1'b0, 10'd342},{8'd129, 1'b1, 10'd349},
{8'd128, 1'b0, 10'd336},{8'd128, 1'b1, 10'd343},
{8'd127, 1'b0, 10'd330},{8'd127, 1'b1, 10'd337},
{8'd126, 1'b0, 10'd324},{8'd126, 1'b1, 10'd331},
{8'd125, 1'b0, 10'd318},{8'd125, 1'b1, 10'd325},
{8'd124, 1'b0, 10'd312},{8'd124, 1'b1, 10'd319},
{8'd123, 1'b0, 10'd306},{8'd123, 1'b1, 10'd313},
{8'd122, 1'b0, 10'd300},{8'd122, 1'b1, 10'd307},
{8'd121, 1'b0, 10'd294},{8'd121, 1'b1, 10'd301},
{8'd120, 1'b0, 10'd288},{8'd120, 1'b1, 10'd295},
{8'd119, 1'b0, 10'd282},{8'd119, 1'b1, 10'd289},
{8'd118, 1'b0, 10'd276},{8'd118, 1'b1, 10'd283},
{8'd117, 1'b0, 10'd270},{8'd117, 1'b1, 10'd277},
{8'd116, 1'b0, 10'd264},{8'd116, 1'b1, 10'd271},
{8'd115, 1'b0, 10'd258},{8'd115, 1'b1, 10'd265},
{8'd114, 1'b0, 10'd252},{8'd114, 1'b1, 10'd259},
{8'd113, 1'b0, 10'd246},{8'd113, 1'b1, 10'd253},
{8'd112, 1'b0, 10'd240},{8'd112, 1'b1, 10'd247},
{8'd111, 1'b0, 10'd234},{8'd111, 1'b1, 10'd241},
{8'd110, 1'b0, 10'd228},{8'd110, 1'b1, 10'd235},
{8'd109, 1'b0, 10'd222},{8'd109, 1'b1, 10'd229},
{8'd108, 1'b0, 10'd216},{8'd108, 1'b1, 10'd223},
{8'd107, 1'b0, 10'd210},{8'd107, 1'b1, 10'd217},
{8'd106, 1'b0, 10'd204},{8'd106, 1'b1, 10'd211},
{8'd105, 1'b0, 10'd198},{8'd105, 1'b1, 10'd205},
{8'd104, 1'b0, 10'd192},{8'd104, 1'b1, 10'd199},
{8'd103, 1'b0, 10'd186},{8'd103, 1'b1, 10'd193},
{8'd102, 1'b0, 10'd180},{8'd102, 1'b1, 10'd187},
{8'd101, 1'b0, 10'd174},{8'd101, 1'b1, 10'd181},
{8'd100, 1'b0, 10'd168},{8'd100, 1'b1, 10'd175},
{ 8'd99, 1'b0, 10'd162},{ 8'd99, 1'b1, 10'd169},
{ 8'd98, 1'b0, 10'd156},{ 8'd98, 1'b1, 10'd163},
{ 8'd97, 1'b0, 10'd150},{ 8'd97, 1'b1, 10'd157},
{ 8'd96, 1'b0, 10'd144},{ 8'd96, 1'b1, 10'd151},
{ 8'd95, 1'b0, 10'd138},{ 8'd95, 1'b1, 10'd145},
{ 8'd94, 1'b0, 10'd132},{ 8'd94, 1'b1, 10'd139},
{ 8'd93, 1'b0, 10'd126},{ 8'd93, 1'b1, 10'd133},
{ 8'd92, 1'b0, 10'd120},{ 8'd92, 1'b1, 10'd127},
{ 8'd91, 1'b0, 10'd114},{ 8'd91, 1'b1, 10'd121},
{ 8'd90, 1'b0, 10'd108},{ 8'd90, 1'b1, 10'd115},
{ 8'd89, 1'b0, 10'd102},{ 8'd89, 1'b1, 10'd109},
{ 8'd88, 1'b0,  10'd96},{ 8'd88, 1'b1, 10'd103},
{ 8'd87, 1'b0,  10'd90},{ 8'd87, 1'b1,  10'd97},
{ 8'd86, 1'b0,  10'd84},{ 8'd86, 1'b1,  10'd91},
{ 8'd85, 1'b0,  10'd78},{ 8'd85, 1'b1,  10'd85},
{ 8'd84, 1'b0,  10'd72},{ 8'd84, 1'b1,  10'd79},
{ 8'd83, 1'b0,  10'd66},{ 8'd83, 1'b1,  10'd73},
{ 8'd82, 1'b0,  10'd60},{ 8'd82, 1'b1,  10'd67},
{ 8'd81, 1'b0,  10'd54},{ 8'd81, 1'b1,  10'd61},
{ 8'd80, 1'b0,  10'd48},{ 8'd80, 1'b1,  10'd55},
{ 8'd79, 1'b0,  10'd42},{ 8'd79, 1'b1,  10'd49},
{ 8'd78, 1'b0,  10'd36},{ 8'd78, 1'b1,  10'd43},
{ 8'd77, 1'b0,  10'd30},{ 8'd77, 1'b1,  10'd37},
{ 8'd76, 1'b0,  10'd24},{ 8'd76, 1'b1,  10'd31},
{ 8'd75, 1'b0,  10'd18},{ 8'd75, 1'b1,  10'd25},
{ 8'd74, 1'b0,  10'd12},{ 8'd74, 1'b1,  10'd19},
{ 8'd73, 1'b0,   10'd6},{ 8'd73, 1'b1,  10'd13},
{ 8'd72, 1'b0,   10'd1},{ 8'd72, 1'b1,   10'd7},
{ 8'd71, 1'b0,   10'd2},{ 8'd71, 1'b0,  10'd26},{ 8'd71, 1'b1, 10'd476},
{ 8'd70, 1'b0, 10'd464},{ 8'd70, 1'b0, 10'd470},{ 8'd70, 1'b1, 10'd560},
{ 8'd69, 1'b0, 10'd200},{ 8'd69, 1'b0, 10'd266},{ 8'd69, 1'b1, 10'd314},
{ 8'd68, 1'b0, 10'd116},{ 8'd68, 1'b0, 10'd260},{ 8'd68, 1'b1, 10'd284},
{ 8'd67, 1'b0,  10'd62},{ 8'd67, 1'b0, 10'd212},{ 8'd67, 1'b1, 10'd500},
{ 8'd66, 1'b0,  10'd32},{ 8'd66, 1'b0, 10'd380},{ 8'd66, 1'b1, 10'd524},
{ 8'd65, 1'b0, 10'd140},{ 8'd65, 1'b0, 10'd224},{ 8'd65, 1'b1, 10'd512},
{ 8'd64, 1'b0, 10'd176},{ 8'd64, 1'b0, 10'd344},{ 8'd64, 1'b1, 10'd632},
{ 8'd63, 1'b0, 10'd110},{ 8'd63, 1'b0, 10'd488},{ 8'd63, 1'b1, 10'd638},
{ 8'd62, 1'b0, 10'd230},{ 8'd62, 1'b0, 10'd320},{ 8'd62, 1'b1, 10'd626},
{ 8'd61, 1'b0,  10'd44},{ 8'd61, 1'b0, 10'd482},{ 8'd61, 1'b1, 10'd590},
{ 8'd60, 1'b0,  10'd80},{ 8'd60, 1'b0, 10'd518},{ 8'd60, 1'b1, 10'd572},
{ 8'd59, 1'b0,  10'd98},{ 8'd59, 1'b0, 10'd104},{ 8'd59, 1'b1, 10'd122},
{ 8'd58, 1'b0, 10'd254},{ 8'd58, 1'b0, 10'd278},{ 8'd58, 1'b1, 10'd398},
{ 8'd57, 1'b0,  10'd92},{ 8'd57, 1'b0, 10'd206},{ 8'd57, 1'b1, 10'd332},
{ 8'd56, 1'b0, 10'd134},{ 8'd56, 1'b0, 10'd152},{ 8'd56, 1'b1, 10'd584},
{ 8'd55, 1'b0, 10'd434},{ 8'd55, 1'b0, 10'd536},{ 8'd55, 1'b1, 10'd542},
{ 8'd54, 1'b0, 10'd428},{ 8'd54, 1'b0, 10'd554},{ 8'd54, 1'b1, 10'd620},
{ 8'd53, 1'b0, 10'd158},{ 8'd53, 1'b0, 10'd188},{ 8'd53, 1'b1, 10'd446},
{ 8'd52, 1'b0, 10'd302},{ 8'd52, 1'b0, 10'd338},{ 8'd52, 1'b1, 10'd506},
{ 8'd51, 1'b0, 10'd182},{ 8'd51, 1'b0, 10'd356},{ 8'd51, 1'b1, 10'd392},
{ 8'd50, 1'b0, 10'd170},{ 8'd50, 1'b0, 10'd242},{ 8'd50, 1'b1, 10'd248},
{ 8'd49, 1'b0,  10'd20},{ 8'd49, 1'b0, 10'd146},{ 8'd49, 1'b1, 10'd416},
{ 8'd48, 1'b0, 10'd128},{ 8'd48, 1'b0, 10'd218},{ 8'd48, 1'b1, 10'd452},
{ 8'd47, 1'b0,  10'd86},{ 8'd47, 1'b0, 10'd350},{ 8'd47, 1'b1, 10'd608},
{ 8'd46, 1'b0,  10'd50},{ 8'd46, 1'b0,  10'd74},{ 8'd46, 1'b1, 10'd368},
{ 8'd45, 1'b0,   10'd8},{ 8'd45, 1'b0, 10'd386},{ 8'd45, 1'b1, 10'd566},
{ 8'd44, 1'b0,  10'd38},{ 8'd44, 1'b0, 10'd308},{ 8'd44, 1'b1, 10'd614},
{ 8'd43, 1'b0,  10'd56},{ 8'd43, 1'b0, 10'd440},{ 8'd43, 1'b1, 10'd578},
{ 8'd42, 1'b0,  10'd68},{ 8'd42, 1'b0, 10'd410},{ 8'd42, 1'b1, 10'd422},
{ 8'd41, 1'b0, 10'd290},{ 8'd41, 1'b0, 10'd362},{ 8'd41, 1'b1, 10'd644},
{ 8'd40, 1'b0,  10'd14},{ 8'd40, 1'b0, 10'd374},{ 8'd40, 1'b1, 10'd596},
{ 8'd39, 1'b0, 10'd164},{ 8'd39, 1'b0, 10'd494},{ 8'd39, 1'b1, 10'd602},
{ 8'd38, 1'b0, 10'd194},{ 8'd38, 1'b0, 10'd326},{ 8'd38, 1'b1, 10'd458},
{ 8'd37, 1'b0, 10'd236},{ 8'd37, 1'b0, 10'd272},{ 8'd37, 1'b1, 10'd296},
{ 8'd36, 1'b0, 10'd404},{ 8'd36, 1'b0, 10'd530},{ 8'd36, 1'b1, 10'd548},
{ 8'd35, 1'b0, 10'd357},{ 8'd35, 1'b0, 10'd417},{ 8'd35, 1'b1, 10'd591},
{ 8'd34, 1'b0, 10'd171},{ 8'd34, 1'b0, 10'd309},{ 8'd34, 1'b1, 10'd633},
{ 8'd33, 1'b0, 10'd225},{ 8'd33, 1'b0, 10'd363},{ 8'd33, 1'b1, 10'd411},
{ 8'd32, 1'b0,   10'd3},{ 8'd32, 1'b0,  10'd45},{ 8'd32, 1'b1, 10'd279},
{ 8'd31, 1'b0, 10'd201},{ 8'd31, 1'b0, 10'd447},{ 8'd31, 1'b1, 10'd465},
{ 8'd30, 1'b0, 10'd405},{ 8'd30, 1'b0, 10'd453},{ 8'd30, 1'b1, 10'd549},
{ 8'd29, 1'b0, 10'd393},{ 8'd29, 1'b0, 10'd454},{ 8'd29, 1'b1, 10'd603},
{ 8'd28, 1'b0,  10'd15},{ 8'd28, 1'b0, 10'd525},{ 8'd28, 1'b1, 10'd579},
{ 8'd27, 1'b0,  10'd87},{ 8'd27, 1'b0, 10'd189},{ 8'd27, 1'b1, 10'd315},
{ 8'd26, 1'b0,  10'd88},{ 8'd26, 1'b0, 10'd531},{ 8'd26, 1'b1, 10'd580},
{ 8'd25, 1'b0, 10'd261},{ 8'd25, 1'b0, 10'd339},{ 8'd25, 1'b1, 10'd555},
{ 8'd24, 1'b0,  10'd46},{ 8'd24, 1'b0, 10'd153},{ 8'd24, 1'b1, 10'd459},
{ 8'd23, 1'b0,   10'd9},{ 8'd23, 1'b0,  10'd21},{ 8'd23, 1'b0,  10'd93},{ 8'd23, 1'b0, 10'd105},{ 8'd23, 1'b0, 10'd177},{ 8'd23, 1'b0, 10'd280},{ 8'd23, 1'b0, 10'd303},{ 8'd23, 1'b0, 10'd375},{ 8'd23, 1'b0, 10'd429},{ 8'd23, 1'b0, 10'd495},{ 8'd23, 1'b0, 10'd537},{ 8'd23, 1'b1, 10'd581},
{ 8'd22, 1'b0,  10'd94},{ 8'd22, 1'b0, 10'd129},{ 8'd22, 1'b0, 10'd165},{ 8'd22, 1'b0, 10'd243},{ 8'd22, 1'b0, 10'd321},{ 8'd22, 1'b0, 10'd345},{ 8'd22, 1'b0, 10'd381},{ 8'd22, 1'b0, 10'd466},{ 8'd22, 1'b0, 10'd489},{ 8'd22, 1'b0, 10'd561},{ 8'd22, 1'b0, 10'd627},{ 8'd22, 1'b1, 10'd634},
{ 8'd21, 1'b0,  10'd63},{ 8'd21, 1'b0,  10'd75},{ 8'd21, 1'b0,  10'd99},{ 8'd21, 1'b0, 10'd111},{ 8'd21, 1'b0, 10'd213},{ 8'd21, 1'b0, 10'd291},{ 8'd21, 1'b0, 10'd435},{ 8'd21, 1'b0, 10'd467},{ 8'd21, 1'b0, 10'd585},{ 8'd21, 1'b0, 10'd609},{ 8'd21, 1'b0, 10'd621},{ 8'd21, 1'b1, 10'd622},
{ 8'd20, 1'b0,  10'd51},{ 8'd20, 1'b0, 10'd297},{ 8'd20, 1'b0, 10'd369},{ 8'd20, 1'b0, 10'd441},{ 8'd20, 1'b0, 10'd496},{ 8'd20, 1'b0, 10'd497},{ 8'd20, 1'b0, 10'd507},{ 8'd20, 1'b0, 10'd508},{ 8'd20, 1'b0, 10'd526},{ 8'd20, 1'b0, 10'd567},{ 8'd20, 1'b0, 10'd586},{ 8'd20, 1'b1, 10'd615},
{ 8'd19, 1'b0,  10'd10},{ 8'd19, 1'b0,  10'd57},{ 8'd19, 1'b0, 10'd154},{ 8'd19, 1'b0, 10'd159},{ 8'd19, 1'b0, 10'd249},{ 8'd19, 1'b0, 10'd285},{ 8'd19, 1'b0, 10'd333},{ 8'd19, 1'b0, 10'd382},{ 8'd19, 1'b0, 10'd387},{ 8'd19, 1'b0, 10'd418},{ 8'd19, 1'b0, 10'd423},{ 8'd19, 1'b1, 10'd490},
{ 8'd18, 1'b0,  10'd64},{ 8'd18, 1'b0, 10'd183},{ 8'd18, 1'b0, 10'd195},{ 8'd18, 1'b0, 10'd255},{ 8'd18, 1'b0, 10'd262},{ 8'd18, 1'b0, 10'd322},{ 8'd18, 1'b0, 10'd334},{ 8'd18, 1'b0, 10'd383},{ 8'd18, 1'b0, 10'd436},{ 8'd18, 1'b0, 10'd455},{ 8'd18, 1'b0, 10'd477},{ 8'd18, 1'b1, 10'd513},
{ 8'd17, 1'b0,  10'd11},{ 8'd17, 1'b0,  10'd39},{ 8'd17, 1'b0,  10'd40},{ 8'd17, 1'b0,  10'd69},{ 8'd17, 1'b0, 10'd100},{ 8'd17, 1'b0, 10'd202},{ 8'd17, 1'b0, 10'd219},{ 8'd17, 1'b0, 10'd323},{ 8'd17, 1'b0, 10'd527},{ 8'd17, 1'b0, 10'd592},{ 8'd17, 1'b0, 10'd597},{ 8'd17, 1'b1, 10'd610},
{ 8'd16, 1'b0,  10'd27},{ 8'd16, 1'b0, 10'd135},{ 8'd16, 1'b0, 10'd155},{ 8'd16, 1'b0, 10'd166},{ 8'd16, 1'b0, 10'd244},{ 8'd16, 1'b0, 10'd267},{ 8'd16, 1'b0, 10'd346},{ 8'd16, 1'b0, 10'd394},{ 8'd16, 1'b0, 10'd399},{ 8'd16, 1'b0, 10'd412},{ 8'd16, 1'b0, 10'd562},{ 8'd16, 1'b1, 10'd598},
{ 8'd15, 1'b0,  10'd70},{ 8'd15, 1'b0, 10'd101},{ 8'd15, 1'b0, 10'd196},{ 8'd15, 1'b0, 10'd207},{ 8'd15, 1'b0, 10'd220},{ 8'd15, 1'b0, 10'd268},{ 8'd15, 1'b0, 10'd460},{ 8'd15, 1'b0, 10'd519},{ 8'd15, 1'b0, 10'd543},{ 8'd15, 1'b0, 10'd604},{ 8'd15, 1'b0, 10'd611},{ 8'd15, 1'b1, 10'd645},
{ 8'd14, 1'b0,  10'd33},{ 8'd14, 1'b0,  10'd89},{ 8'd14, 1'b0,  10'd95},{ 8'd14, 1'b0, 10'd130},{ 8'd14, 1'b0, 10'd286},{ 8'd14, 1'b0, 10'd370},{ 8'd14, 1'b0, 10'd471},{ 8'd14, 1'b0, 10'd520},{ 8'd14, 1'b0, 10'd550},{ 8'd14, 1'b0, 10'd573},{ 8'd14, 1'b0, 10'd599},{ 8'd14, 1'b1, 10'd616},
{ 8'd13, 1'b0,  10'd28},{ 8'd13, 1'b0, 10'd123},{ 8'd13, 1'b0, 10'd214},{ 8'd13, 1'b0, 10'd231},{ 8'd13, 1'b0, 10'd237},{ 8'd13, 1'b0, 10'd256},{ 8'd13, 1'b0, 10'd273},{ 8'd13, 1'b0, 10'd310},{ 8'd13, 1'b0, 10'd327},{ 8'd13, 1'b0, 10'd472},{ 8'd13, 1'b0, 10'd568},{ 8'd13, 1'b1, 10'd623},
{ 8'd12, 1'b0,  10'd22},{ 8'd12, 1'b0,  10'd52},{ 8'd12, 1'b0,  10'd71},{ 8'd12, 1'b0, 10'd136},{ 8'd12, 1'b0, 10'd232},{ 8'd12, 1'b0, 10'd316},{ 8'd12, 1'b0, 10'd347},{ 8'd12, 1'b0, 10'd358},{ 8'd12, 1'b0, 10'd400},{ 8'd12, 1'b0, 10'd448},{ 8'd12, 1'b0, 10'd449},{ 8'd12, 1'b1, 10'd478},
{ 8'd11, 1'b0,  10'd16},{ 8'd11, 1'b0,  10'd65},{ 8'd11, 1'b0, 10'd117},{ 8'd11, 1'b0, 10'd190},{ 8'd11, 1'b0, 10'd226},{ 8'd11, 1'b0, 10'd238},{ 8'd11, 1'b0, 10'd263},{ 8'd11, 1'b0, 10'd274},{ 8'd11, 1'b0, 10'd298},{ 8'd11, 1'b0, 10'd364},{ 8'd11, 1'b0, 10'd371},{ 8'd11, 1'b1, 10'd430},
{ 8'd10, 1'b0,  10'd41},{ 8'd10, 1'b0,  10'd58},{ 8'd10, 1'b0, 10'd141},{ 8'd10, 1'b0, 10'd208},{ 8'd10, 1'b0, 10'd351},{ 8'd10, 1'b0, 10'd473},{ 8'd10, 1'b0, 10'd491},{ 8'd10, 1'b0, 10'd501},{ 8'd10, 1'b0, 10'd514},{ 8'd10, 1'b0, 10'd521},{ 8'd10, 1'b0, 10'd538},{ 8'd10, 1'b1, 10'd574},
{  8'd9, 1'b0,  10'd47},{  8'd9, 1'b0, 10'd112},{  8'd9, 1'b0, 10'd142},{  8'd9, 1'b0, 10'd197},{  8'd9, 1'b0, 10'd203},{  8'd9, 1'b0, 10'd221},{  8'd9, 1'b0, 10'd317},{  8'd9, 1'b0, 10'd328},{  8'd9, 1'b0, 10'd359},{  8'd9, 1'b0, 10'd532},{  8'd9, 1'b0, 10'd556},{  8'd9, 1'b1, 10'd639},
{  8'd8, 1'b0,  10'd53},{  8'd8, 1'b0,  10'd81},{  8'd8, 1'b0, 10'd106},{  8'd8, 1'b0, 10'd118},{  8'd8, 1'b0, 10'd160},{  8'd8, 1'b0, 10'd172},{  8'd8, 1'b0, 10'd233},{  8'd8, 1'b0, 10'd335},{  8'd8, 1'b0, 10'd340},{  8'd8, 1'b0, 10'd406},{  8'd8, 1'b0, 10'd424},{  8'd8, 1'b1, 10'd442},
{  8'd7, 1'b0,  10'd82},{  8'd7, 1'b0, 10'd113},{  8'd7, 1'b0, 10'd131},{  8'd7, 1'b0, 10'd245},{  8'd7, 1'b0, 10'd269},{  8'd7, 1'b0, 10'd341},{  8'd7, 1'b0, 10'd419},{  8'd7, 1'b0, 10'd483},{  8'd7, 1'b0, 10'd484},{  8'd7, 1'b0, 10'd593},{  8'd7, 1'b0, 10'd628},{  8'd7, 1'b1, 10'd646},
{  8'd6, 1'b0,  10'd17},{  8'd6, 1'b0, 10'd119},{  8'd6, 1'b0, 10'd173},{  8'd6, 1'b0, 10'd184},{  8'd6, 1'b0, 10'd191},{  8'd6, 1'b0, 10'd215},{  8'd6, 1'b0, 10'd287},{  8'd6, 1'b0, 10'd329},{  8'd6, 1'b0, 10'd376},{  8'd6, 1'b0, 10'd515},{  8'd6, 1'b0, 10'd539},{  8'd6, 1'b1, 10'd544},
{  8'd5, 1'b0,  10'd29},{  8'd5, 1'b0,  10'd34},{  8'd5, 1'b0, 10'd124},{  8'd5, 1'b0, 10'd147},{  8'd5, 1'b0, 10'd250},{  8'd5, 1'b0, 10'd365},{  8'd5, 1'b0, 10'd388},{  8'd5, 1'b0, 10'd395},{  8'd5, 1'b0, 10'd502},{  8'd5, 1'b0, 10'd557},{  8'd5, 1'b0, 10'd617},{  8'd5, 1'b1, 10'd640},
{  8'd4, 1'b0,  10'd35},{  8'd4, 1'b0, 10'd107},{  8'd4, 1'b0, 10'd148},{  8'd4, 1'b0, 10'd161},{  8'd4, 1'b0, 10'd178},{  8'd4, 1'b0, 10'd239},{  8'd4, 1'b0, 10'd251},{  8'd4, 1'b0, 10'd377},{  8'd4, 1'b0, 10'd389},{  8'd4, 1'b0, 10'd413},{  8'd4, 1'b0, 10'd533},{  8'd4, 1'b1, 10'd605},
{  8'd3, 1'b0, 10'd149},{  8'd3, 1'b0, 10'd185},{  8'd3, 1'b0, 10'd299},{  8'd3, 1'b0, 10'd304},{  8'd3, 1'b0, 10'd311},{  8'd3, 1'b0, 10'd401},{  8'd3, 1'b0, 10'd461},{  8'd3, 1'b0, 10'd479},{  8'd3, 1'b0, 10'd545},{  8'd3, 1'b0, 10'd551},{  8'd3, 1'b0, 10'd587},{  8'd3, 1'b1, 10'd635},
{  8'd2, 1'b0,  10'd59},{  8'd2, 1'b0,  10'd76},{  8'd2, 1'b0, 10'd137},{  8'd2, 1'b0, 10'd227},{  8'd2, 1'b0, 10'd275},{  8'd2, 1'b0, 10'd292},{  8'd2, 1'b0, 10'd352},{  8'd2, 1'b0, 10'd353},{  8'd2, 1'b0, 10'd437},{  8'd2, 1'b0, 10'd485},{  8'd2, 1'b0, 10'd575},{  8'd2, 1'b1, 10'd647},
{  8'd1, 1'b0,  10'd23},{  8'd1, 1'b0, 10'd125},{  8'd1, 1'b0, 10'd167},{  8'd1, 1'b0, 10'd179},{  8'd1, 1'b0, 10'd305},{  8'd1, 1'b0, 10'd407},{  8'd1, 1'b0, 10'd425},{  8'd1, 1'b0, 10'd443},{  8'd1, 1'b0, 10'd509},{  8'd1, 1'b0, 10'd569},{  8'd1, 1'b0, 10'd629},{  8'd1, 1'b1, 10'd641},
{  8'd0, 1'b0,   10'd4},{  8'd0, 1'b0,   10'd5},{  8'd0, 1'b0,  10'd77},{  8'd0, 1'b0,  10'd83},{  8'd0, 1'b0, 10'd143},{  8'd0, 1'b0, 10'd209},{  8'd0, 1'b0, 10'd257},{  8'd0, 1'b0, 10'd281},{  8'd0, 1'b0, 10'd293},{  8'd0, 1'b0, 10'd431},{  8'd0, 1'b0, 10'd503},{  8'd0, 1'b1, 10'd563}
};
localparam int          cLARGE_HS_TAB_1BY2_PACKED_SIZE = 630;
localparam bit [18 : 0] cLARGE_HS_TAB_1BY2_PACKED[cLARGE_HS_TAB_1BY2_PACKED_SIZE] = '{
{  1'b1, 1'b0, 8'd179,    9'd1},{  1'b0, 1'b0,  8'd90,    9'd0},{  1'b0, 1'b0,  8'd74,  9'd181},{  1'b0, 1'b0,  8'd36,    9'd0},{  1'b0, 1'b0,  8'd30,   9'd67},{  1'b0, 1'b0,  8'd27,  9'd259},{  1'b0, 1'b1,  8'd26,  9'd300},
{  1'b0, 1'b0,  8'd91,    9'd0},{  1'b0, 1'b0,  8'd90,    9'd0},{  1'b0, 1'b0,  8'd41,  9'd154},{  1'b0, 1'b0,  8'd37,    9'd0},{  1'b0, 1'b0,  8'd20,  9'd286},{  1'b0, 1'b0,  8'd10,   9'd50},{  1'b0, 1'b1,  8'd10,   9'd61},
{  1'b0, 1'b0,  8'd92,    9'd0},{  1'b0, 1'b0,  8'd91,    9'd0},{  1'b0, 1'b0,  8'd51,  9'd138},{  1'b0, 1'b0,  8'd38,    9'd0},{  1'b0, 1'b0,  8'd27,  9'd318},{  1'b0, 1'b0,  8'd16,   9'd14},{  1'b0, 1'b1,   8'd4,   9'd31},
{  1'b0, 1'b0,  8'd93,    9'd0},{  1'b0, 1'b0,  8'd92,    9'd0},{  1'b0, 1'b0,  8'd68,  9'd352},{  1'b0, 1'b0,  8'd39,    9'd0},{  1'b0, 1'b0,  8'd16,  9'd267},{  1'b0, 1'b0,   8'd6,   9'd69},{  1'b0, 1'b1,   8'd2,  9'd262},
{  1'b0, 1'b0,  8'd94,    9'd0},{  1'b0, 1'b0,  8'd93,    9'd0},{  1'b0, 1'b0,  8'd82,  9'd278},{  1'b0, 1'b0,  8'd40,    9'd0},{  1'b0, 1'b0,  8'd33,   9'd36},{  1'b0, 1'b0,  8'd24,  9'd239},{  1'b0, 1'b1,   8'd9,  9'd317},
{  1'b0, 1'b0,  8'd95,    9'd0},{  1'b0, 1'b0,  8'd94,    9'd0},{  1'b0, 1'b0,  8'd41,    9'd0},{  1'b0, 1'b0,  8'd30,  9'd209},{  1'b0, 1'b0,  8'd24,  9'd136},{  1'b0, 1'b0,  8'd13,  9'd254},{  1'b0, 1'b1,   8'd3,  9'd152},
{  1'b0, 1'b0,  8'd96,    9'd0},{  1'b0, 1'b0,  8'd95,    9'd0},{  1'b0, 1'b0,  8'd76,  9'd338},{  1'b0, 1'b0,  8'd42,    9'd0},{  1'b0, 1'b0,  8'd32,  9'd236},{  1'b0, 1'b0,  8'd21,  9'd103},{  1'b0, 1'b1,  8'd14,  9'd286},
{  1'b0, 1'b0,  8'd97,    9'd0},{  1'b0, 1'b0,  8'd96,    9'd0},{  1'b0, 1'b0,  8'd89,  9'd214},{  1'b0, 1'b0,  8'd43,    9'd0},{  1'b0, 1'b0,  8'd34,  9'd265},{  1'b0, 1'b0,  8'd28,   9'd44},{  1'b0, 1'b1,   8'd4,  9'd126},
{  1'b0, 1'b0,  8'd98,    9'd0},{  1'b0, 1'b0,  8'd97,    9'd0},{  1'b0, 1'b0,  8'd87,   9'd49},{  1'b0, 1'b0,  8'd44,    9'd0},{  1'b0, 1'b0,  8'd30,  9'd297},{  1'b0, 1'b0,  8'd18,   9'd15},{  1'b0, 1'b1,  8'd16,  9'd332},
{  1'b0, 1'b0,  8'd99,    9'd0},{  1'b0, 1'b0,  8'd98,    9'd0},{  1'b0, 1'b0,  8'd79,  9'd353},{  1'b0, 1'b0,  8'd58,  9'd296},{  1'b0, 1'b0,  8'd45,    9'd0},{  1'b0, 1'b0,  8'd24,  9'd341},{  1'b0, 1'b1,  8'd21,  9'd341},
{  1'b0, 1'b0, 8'd100,    9'd0},{  1'b0, 1'b0,  8'd99,    9'd0},{  1'b0, 1'b0,  8'd46,    9'd0},{  1'b0, 1'b0,  8'd37,    9'd1},{  1'b0, 1'b0,   8'd5,  9'd176},{  1'b0, 1'b0,   8'd4,  9'd140},{  1'b0, 1'b1,   8'd1,   9'd28},
{  1'b0, 1'b0, 8'd101,    9'd0},{  1'b0, 1'b0, 8'd100,    9'd0},{  1'b0, 1'b0,  8'd47,    9'd0},{  1'b0, 1'b0,  8'd32,  9'd170},{  1'b0, 1'b0,  8'd20,  9'd133},{  1'b0, 1'b0,  8'd19,  9'd200},{  1'b0, 1'b1,   8'd8,  9'd277},
{  1'b0, 1'b0, 8'd102,    9'd0},{  1'b0, 1'b0, 8'd101,    9'd0},{  1'b0, 1'b0,  8'd78,  9'd197},{  1'b0, 1'b0,  8'd48,    9'd0},{  1'b0, 1'b0,  8'd33,  9'd181},{  1'b0, 1'b0,  8'd26,   9'd79},{  1'b0, 1'b1,  8'd15,  9'd333},
{  1'b0, 1'b0, 8'd103,    9'd0},{  1'b0, 1'b0, 8'd102,    9'd0},{  1'b0, 1'b0,  8'd66,  9'd231},{  1'b0, 1'b0,  8'd49,    9'd0},{  1'b0, 1'b0,  8'd46,  9'd315},{  1'b0, 1'b0,  8'd16,  9'd145},{  1'b0, 1'b1,   8'd8,  9'd100},
{  1'b0, 1'b0, 8'd104,    9'd0},{  1'b0, 1'b0, 8'd103,    9'd0},{  1'b0, 1'b0,  8'd67,  9'd131},{  1'b0, 1'b0,  8'd63,  9'd100},{  1'b0, 1'b0,  8'd50,    9'd0},{  1'b0, 1'b0,  8'd18,  9'd226},{  1'b0, 1'b1,   8'd0,   9'd28},
{  1'b0, 1'b0, 8'd105,    9'd0},{  1'b0, 1'b0, 8'd104,    9'd0},{  1'b0, 1'b0,  8'd63,  9'd299},{  1'b0, 1'b0,  8'd51,    9'd0},{  1'b0, 1'b0,  8'd30,  9'd184},{  1'b0, 1'b0,  8'd23,  9'd335},{  1'b0, 1'b1,  8'd13,  9'd166},
{  1'b0, 1'b0, 8'd106,    9'd0},{  1'b0, 1'b0, 8'd105,    9'd0},{  1'b0, 1'b0,  8'd73,   9'd85},{  1'b0, 1'b0,  8'd59,  9'd124},{  1'b0, 1'b0,  8'd52,    9'd0},{  1'b0, 1'b0,  8'd11,  9'd239},{  1'b0, 1'b1,   8'd6,  9'd135},
{  1'b0, 1'b0, 8'd107,    9'd0},{  1'b0, 1'b0, 8'd106,    9'd0},{  1'b0, 1'b0,  8'd56,  9'd302},{  1'b0, 1'b0,  8'd53,    9'd0},{  1'b0, 1'b0,  8'd49,  9'd121},{  1'b0, 1'b0,  8'd27,   9'd54},{  1'b0, 1'b1,   8'd8,  9'd173},
{  1'b0, 1'b0, 8'd108,    9'd0},{  1'b0, 1'b0, 8'd107,    9'd0},{  1'b0, 1'b0,  8'd81,  9'd161},{  1'b0, 1'b0,  8'd54,    9'd0},{  1'b0, 1'b0,  8'd25,  9'd273},{  1'b0, 1'b0,  8'd23,   9'd51},{  1'b0, 1'b1,  8'd14,  9'd110},
{  1'b0, 1'b0, 8'd109,    9'd0},{  1'b0, 1'b0, 8'd108,    9'd0},{  1'b0, 1'b0,  8'd55,    9'd0},{  1'b0, 1'b0,  8'd38,  9'd114},{  1'b0, 1'b0,  8'd28,  9'd160},{  1'b0, 1'b0,  8'd15,  9'd139},{  1'b0, 1'b1,   8'd2,  9'd192},
{  1'b0, 1'b0, 8'd110,    9'd0},{  1'b0, 1'b0, 8'd109,    9'd0},{  1'b0, 1'b0,  8'd74,   9'd94},{  1'b0, 1'b0,  8'd56,    9'd0},{  1'b0, 1'b0,  8'd31,  9'd293},{  1'b0, 1'b0,  8'd19,   9'd34},{  1'b0, 1'b1,  8'd11,   9'd50},
{  1'b0, 1'b0, 8'd111,    9'd0},{  1'b0, 1'b0, 8'd110,    9'd0},{  1'b0, 1'b0,  8'd67,  9'd280},{  1'b0, 1'b0,  8'd57,    9'd0},{  1'b0, 1'b0,  8'd11,  9'd188},{  1'b0, 1'b0,   8'd8,   9'd23},{  1'b0, 1'b1,   8'd0,  9'd306},
{  1'b0, 1'b0, 8'd112,    9'd0},{  1'b0, 1'b0, 8'd111,    9'd0},{  1'b0, 1'b0,  8'd85,   9'd55},{  1'b0, 1'b0,  8'd71,  9'd290},{  1'b0, 1'b0,  8'd58,    9'd0},{  1'b0, 1'b0,  8'd31,  9'd306},{  1'b0, 1'b1,  8'd19,   9'd89},
{  1'b0, 1'b0, 8'd113,    9'd0},{  1'b0, 1'b0, 8'd112,    9'd0},{  1'b0, 1'b0,  8'd59,    9'd0},{  1'b0, 1'b0,  8'd45,  9'd184},{  1'b0, 1'b0,  8'd19,  9'd170},{  1'b0, 1'b0,   8'd9,   9'd44},{  1'b0, 1'b1,   8'd3,  9'd207},
{  1'b0, 1'b0, 8'd114,    9'd0},{  1'b0, 1'b0, 8'd113,    9'd0},{  1'b0, 1'b0,  8'd60,    9'd0},{  1'b0, 1'b0,  8'd52,   9'd97},{  1'b0, 1'b0,  8'd35,  9'd204},{  1'b0, 1'b0,  8'd17,   9'd73},{  1'b0, 1'b1,   8'd4,   9'd35},
{  1'b0, 1'b0, 8'd115,    9'd0},{  1'b0, 1'b0, 8'd114,    9'd0},{  1'b0, 1'b0,  8'd78,   9'd76},{  1'b0, 1'b0,  8'd61,    9'd0},{  1'b0, 1'b0,  8'd27,  9'd228},{  1'b0, 1'b0,  8'd24,  9'd289},{  1'b0, 1'b1,  8'd19,    9'd3},
{  1'b0, 1'b0, 8'd116,    9'd0},{  1'b0, 1'b0, 8'd115,    9'd0},{  1'b0, 1'b0,  8'd83,  9'd243},{  1'b0, 1'b0,  8'd62,    9'd0},{  1'b0, 1'b0,  8'd52,   9'd85},{  1'b0, 1'b0,  8'd29,  9'd117},{  1'b0, 1'b1,   8'd2,  9'd289},
{  1'b0, 1'b0, 8'd117,    9'd0},{  1'b0, 1'b0, 8'd116,    9'd0},{  1'b0, 1'b0,  8'd66,   9'd19},{  1'b0, 1'b0,  8'd63,    9'd0},{  1'b0, 1'b0,  8'd34,   9'd69},{  1'b0, 1'b0,  8'd13,  9'd168},{  1'b0, 1'b1,   8'd7,  9'd130},
{  1'b0, 1'b0, 8'd118,    9'd0},{  1'b0, 1'b0, 8'd117,    9'd0},{  1'b0, 1'b0,  8'd64,    9'd0},{  1'b0, 1'b0,  8'd45,  9'd123},{  1'b0, 1'b0,  8'd32,   9'd10},{  1'b0, 1'b0,  8'd25,  9'd332},{  1'b0, 1'b1,  8'd18,  9'd273},
{  1'b0, 1'b0, 8'd119,    9'd0},{  1'b0, 1'b0, 8'd118,    9'd0},{  1'b0, 1'b0,  8'd65,    9'd0},{  1'b0, 1'b0,  8'd35,  9'd141},{  1'b0, 1'b0,  8'd14,   9'd74},{  1'b0, 1'b0,   8'd6,  9'd238},{  1'b0, 1'b1,   8'd5,  9'd238},
{  1'b0, 1'b0, 8'd120,    9'd0},{  1'b0, 1'b0, 8'd119,    9'd0},{  1'b0, 1'b0,  8'd86,   9'd30},{  1'b0, 1'b0,  8'd66,    9'd0},{  1'b0, 1'b0,  8'd47,  9'd155},{  1'b0, 1'b0,  8'd22,   9'd61},{  1'b0, 1'b1,  8'd20,  9'd126},
{  1'b0, 1'b0, 8'd121,    9'd0},{  1'b0, 1'b0, 8'd120,    9'd0},{  1'b0, 1'b0,  8'd80,  9'd233},{  1'b0, 1'b0,  8'd67,    9'd0},{  1'b0, 1'b0,  8'd46,  9'd185},{  1'b0, 1'b0,   8'd4,  9'd326},{  1'b0, 1'b1,   8'd3,  9'd128},
{  1'b0, 1'b0, 8'd122,    9'd0},{  1'b0, 1'b0, 8'd121,    9'd0},{  1'b0, 1'b0,  8'd68,    9'd0},{  1'b0, 1'b0,  8'd64,  9'd213},{  1'b0, 1'b0,  8'd25,  9'd189},{  1'b0, 1'b0,  8'd17,  9'd329},{  1'b0, 1'b1,   8'd6,  9'd202},
{  1'b0, 1'b0, 8'd123,    9'd0},{  1'b0, 1'b0, 8'd122,    9'd0},{  1'b0, 1'b0,  8'd69,    9'd0},{  1'b0, 1'b0,  8'd40,   9'd46},{  1'b0, 1'b0,  8'd35,  9'd293},{  1'b0, 1'b0,  8'd16,   9'd87},{  1'b0, 1'b1,  8'd15,  9'd111},
{  1'b0, 1'b0, 8'd124,    9'd0},{  1'b0, 1'b0, 8'd123,    9'd0},{  1'b0, 1'b0,  8'd88,  9'd324},{  1'b0, 1'b0,  8'd77,  9'd171},{  1'b0, 1'b0,  8'd70,    9'd0},{  1'b0, 1'b0,  8'd12,  9'd288},{  1'b0, 1'b1,  8'd11,   9'd47},
{  1'b0, 1'b0, 8'd125,    9'd0},{  1'b0, 1'b0, 8'd124,    9'd0},{  1'b0, 1'b0,  8'd71,    9'd0},{  1'b0, 1'b0,  8'd36,  9'd277},{  1'b0, 1'b0,  8'd28,  9'd173},{  1'b0, 1'b0,  8'd22,  9'd152},{  1'b0, 1'b1,  8'd14,  9'd229},
{  1'b0, 1'b0, 8'd126,    9'd0},{  1'b0, 1'b0, 8'd125,    9'd0},{  1'b0, 1'b0,  8'd72,    9'd0},{  1'b0, 1'b0,  8'd51,  9'd296},{  1'b0, 1'b0,  8'd25,  9'd277},{  1'b0, 1'b0,  8'd21,  9'd229},{  1'b0, 1'b1,   8'd5,   9'd35},
{  1'b0, 1'b0, 8'd127,    9'd0},{  1'b0, 1'b0, 8'd126,    9'd0},{  1'b0, 1'b0,  8'd73,    9'd0},{  1'b0, 1'b0,  8'd61,  9'd196},{  1'b0, 1'b0,  8'd31,   9'd69},{  1'b0, 1'b0,  8'd10,  9'd285},{  1'b0, 1'b1,   8'd4,  9'd144},
{  1'b0, 1'b0, 8'd128,    9'd0},{  1'b0, 1'b0, 8'd127,    9'd0},{  1'b0, 1'b0,  8'd74,    9'd0},{  1'b0, 1'b0,  8'd50,   9'd42},{  1'b0, 1'b0,  8'd37,   9'd43},{  1'b0, 1'b0,  8'd10,  9'd164},{  1'b0, 1'b1,   8'd7,  9'd103},
{  1'b0, 1'b0, 8'd129,    9'd0},{  1'b0, 1'b0, 8'd128,    9'd0},{  1'b0, 1'b0,  8'd75,    9'd0},{  1'b0, 1'b0,  8'd55,   9'd95},{  1'b0, 1'b0,  8'd48,  9'd357},{  1'b0, 1'b0,  8'd26,  9'd332},{  1'b0, 1'b1,  8'd20,  9'd101},
{  1'b0, 1'b0, 8'd130,    9'd0},{  1'b0, 1'b0, 8'd129,    9'd0},{  1'b0, 1'b0,  8'd76,    9'd0},{  1'b0, 1'b0,  8'd75,  9'd112},{  1'b0, 1'b0,  8'd70,  9'd136},{  1'b0, 1'b0,  8'd20,   9'd88},{  1'b0, 1'b1,  8'd15,  9'd337},
{  1'b0, 1'b0, 8'd131,    9'd0},{  1'b0, 1'b0, 8'd130,    9'd0},{  1'b0, 1'b0,  8'd77,    9'd0},{  1'b0, 1'b0,  8'd58,   9'd67},{  1'b0, 1'b0,  8'd57,  9'd167},{  1'b0, 1'b0,  8'd31,  9'd275},{  1'b0, 1'b1,  8'd17,  9'd349},
{  1'b0, 1'b0, 8'd132,    9'd0},{  1'b0, 1'b0, 8'd131,    9'd0},{  1'b0, 1'b0,  8'd86,   9'd73},{  1'b0, 1'b0,  8'd78,    9'd0},{  1'b0, 1'b0,  8'd27,  9'd245},{  1'b0, 1'b0,  8'd20,  9'd238},{  1'b0, 1'b1,  8'd16,  9'd311},
{  1'b0, 1'b0, 8'd133,    9'd0},{  1'b0, 1'b0, 8'd132,    9'd0},{  1'b0, 1'b0,  8'd89,  9'd223},{  1'b0, 1'b0,  8'd79,    9'd0},{  1'b0, 1'b0,  8'd59,  9'd115},{  1'b0, 1'b0,  8'd21,   9'd50},{  1'b0, 1'b1,  8'd14,   9'd60},
{  1'b0, 1'b0, 8'd134,    9'd0},{  1'b0, 1'b0, 8'd133,    9'd0},{  1'b0, 1'b0,  8'd80,    9'd0},{  1'b0, 1'b0,  8'd39,    9'd8},{  1'b0, 1'b0,  8'd25,  9'd107},{  1'b0, 1'b0,  8'd19,  9'd148},{  1'b0, 1'b1,   8'd8,   9'd60},
{  1'b0, 1'b0, 8'd135,    9'd0},{  1'b0, 1'b0, 8'd134,    9'd0},{  1'b0, 1'b0,  8'd81,    9'd0},{  1'b0, 1'b0,  8'd22,  9'd177},{  1'b0, 1'b0,  8'd18,   9'd58},{  1'b0, 1'b0,   8'd5,   9'd68},{  1'b0, 1'b1,   8'd1,   9'd51},
{  1'b0, 1'b0, 8'd136,    9'd0},{  1'b0, 1'b0, 8'd135,    9'd0},{  1'b0, 1'b0,  8'd82,    9'd0},{  1'b0, 1'b0,  8'd71,   9'd72},{  1'b0, 1'b0,  8'd33,   9'd25},{  1'b0, 1'b0,  8'd21,  9'd329},{  1'b0, 1'b1,   8'd7,   9'd65},
{  1'b0, 1'b0, 8'd137,    9'd0},{  1'b0, 1'b0, 8'd136,    9'd0},{  1'b0, 1'b0,  8'd83,    9'd0},{  1'b0, 1'b0,  8'd65,  9'd340},{  1'b0, 1'b0,  8'd50,  9'd239},{  1'b0, 1'b0,  8'd26,  9'd165},{  1'b0, 1'b1,   8'd0,   9'd95},
{  1'b0, 1'b0, 8'd138,    9'd0},{  1'b0, 1'b0, 8'd137,    9'd0},{  1'b0, 1'b0,  8'd84,    9'd0},{  1'b0, 1'b0,  8'd35,  9'd211},{  1'b0, 1'b0,  8'd14,  9'd204},{  1'b0, 1'b0,  8'd10,  9'd179},{  1'b0, 1'b1,   8'd0,  9'd103},
{  1'b0, 1'b0, 8'd139,    9'd0},{  1'b0, 1'b0, 8'd138,    9'd0},{  1'b0, 1'b0,  8'd85,    9'd0},{  1'b0, 1'b0,  8'd33,  9'd296},{  1'b0, 1'b0,  8'd29,   9'd19},{  1'b0, 1'b0,   8'd5,  9'd186},{  1'b0, 1'b1,   8'd0,  9'd113},
{  1'b0, 1'b0, 8'd140,    9'd0},{  1'b0, 1'b0, 8'd139,    9'd0},{  1'b0, 1'b0,  8'd86,    9'd0},{  1'b0, 1'b0,  8'd60,  9'd148},{  1'b0, 1'b0,  8'd12,  9'd116},{  1'b0, 1'b0,  8'd11,  9'd248},{  1'b0, 1'b1,   8'd1,  9'd312},
{  1'b0, 1'b0, 8'd141,    9'd0},{  1'b0, 1'b0, 8'd140,    9'd0},{  1'b0, 1'b0,  8'd87,    9'd0},{  1'b0, 1'b0,  8'd85,  9'd229},{  1'b0, 1'b0,  8'd21,  9'd243},{  1'b0, 1'b0,   8'd3,   9'd64},{  1'b0, 1'b1,   8'd1,   9'd40},
{  1'b0, 1'b0, 8'd142,    9'd0},{  1'b0, 1'b0, 8'd141,    9'd0},{  1'b0, 1'b0,  8'd88,    9'd0},{  1'b0, 1'b0,  8'd87,  9'd141},{  1'b0, 1'b0,  8'd73,  9'd299},{  1'b0, 1'b0,  8'd17,  9'd350},{  1'b0, 1'b1,   8'd5,  9'd235},
{  1'b0, 1'b0, 8'd143,    9'd0},{  1'b0, 1'b0, 8'd142,    9'd0},{  1'b0, 1'b0,  8'd89,    9'd0},{  1'b0, 1'b0,  8'd68,  9'd197},{  1'b0, 1'b0,  8'd40,  9'd137},{  1'b0, 1'b0,  8'd23,  9'd145},{  1'b0, 1'b1,  8'd10,  9'd246},
{  1'b0, 1'b0, 8'd144,    9'd0},{  1'b0, 1'b0, 8'd143,    9'd0},{  1'b0, 1'b0,  8'd83,   9'd50},{  1'b0, 1'b0,   8'd8,  9'd262},{  1'b0, 1'b0,   8'd6,   9'd92},{  1'b0, 1'b0,   8'd3,  9'd290},{  1'b0, 1'b1,   8'd0,    9'd0},
{  1'b0, 1'b0, 8'd145,    9'd0},{  1'b0, 1'b0, 8'd144,    9'd0},{  1'b0, 1'b0,  8'd88,    9'd6},{  1'b0, 1'b0,  8'd53,  9'd165},{  1'b0, 1'b0,  8'd30,    9'd5},{  1'b0, 1'b0,  8'd25,  9'd347},{  1'b0, 1'b1,   8'd1,    9'd0},
{  1'b0, 1'b0, 8'd146,    9'd0},{  1'b0, 1'b0, 8'd145,    9'd0},{  1'b0, 1'b0,  8'd42,   9'd11},{  1'b0, 1'b0,  8'd30,   9'd32},{  1'b0, 1'b0,  8'd28,  9'd176},{  1'b0, 1'b0,   8'd6,  9'd344},{  1'b0, 1'b1,   8'd2,    9'd0},
{  1'b0, 1'b0, 8'd147,    9'd0},{  1'b0, 1'b0, 8'd146,    9'd0},{  1'b0, 1'b0,  8'd60,  9'd106},{  1'b0, 1'b0,  8'd26,  9'd308},{  1'b0, 1'b0,  8'd12,  9'd106},{  1'b0, 1'b0,   8'd3,    9'd0},{  1'b0, 1'b1,   8'd3,  9'd171},
{  1'b0, 1'b0, 8'd148,    9'd0},{  1'b0, 1'b0, 8'd147,    9'd0},{  1'b0, 1'b0,  8'd35,  9'd279},{  1'b0, 1'b0,  8'd29,   9'd56},{  1'b0, 1'b0,  8'd23,  9'd207},{  1'b0, 1'b0,   8'd4,    9'd0},{  1'b0, 1'b1,   8'd4,  9'd319},
{  1'b0, 1'b0, 8'd149,    9'd0},{  1'b0, 1'b0, 8'd148,    9'd0},{  1'b0, 1'b0,  8'd54,  9'd174},{  1'b0, 1'b0,  8'd44,   9'd89},{  1'b0, 1'b0,  8'd29,  9'd112},{  1'b0, 1'b0,  8'd17,  9'd105},{  1'b0, 1'b1,   8'd5,    9'd0},
{  1'b0, 1'b0, 8'd150,    9'd0},{  1'b0, 1'b0, 8'd149,    9'd0},{  1'b0, 1'b0,  8'd57,  9'd300},{  1'b0, 1'b0,  8'd38,    9'd2},{  1'b0, 1'b0,  8'd21,  9'd311},{  1'b0, 1'b0,  8'd12,  9'd359},{  1'b0, 1'b1,   8'd6,    9'd0},
{  1'b0, 1'b0, 8'd151,    9'd0},{  1'b0, 1'b0, 8'd150,    9'd0},{  1'b0, 1'b0,  8'd70,  9'd295},{  1'b0, 1'b0,  8'd61,   9'd78},{  1'b0, 1'b0,  8'd31,  9'd223},{  1'b0, 1'b0,  8'd12,  9'd342},{  1'b0, 1'b1,   8'd7,    9'd0},
{  1'b0, 1'b0, 8'd152,    9'd0},{  1'b0, 1'b0, 8'd151,    9'd0},{  1'b0, 1'b0,  8'd65,  9'd201},{  1'b0, 1'b0,  8'd35,   9'd98},{  1'b0, 1'b0,  8'd12,   9'd68},{  1'b0, 1'b0,  8'd12,   9'd30},{  1'b0, 1'b1,   8'd8,    9'd0},
{  1'b0, 1'b0, 8'd153,    9'd0},{  1'b0, 1'b0, 8'd152,    9'd0},{  1'b0, 1'b0,  8'd34,  9'd132},{  1'b0, 1'b0,  8'd29,  9'd324},{  1'b0, 1'b0,   8'd9,    9'd0},{  1'b0, 1'b0,   8'd1,   9'd80},{  1'b0, 1'b1,   8'd1,   9'd33},
{  1'b0, 1'b0, 8'd154,    9'd0},{  1'b0, 1'b0, 8'd153,    9'd0},{  1'b0, 1'b0,  8'd33,  9'd225},{  1'b0, 1'b0,  8'd23,  9'd324},{  1'b0, 1'b0,  8'd18,   9'd71},{  1'b0, 1'b0,  8'd10,    9'd0},{  1'b0, 1'b1,   8'd3,  9'd180},
{  1'b0, 1'b0, 8'd155,    9'd0},{  1'b0, 1'b0, 8'd154,    9'd0},{  1'b0, 1'b0,  8'd72,  9'd290},{  1'b0, 1'b0,  8'd47,  9'd274},{  1'b0, 1'b0,  8'd17,  9'd103},{  1'b0, 1'b0,  8'd13,  9'd213},{  1'b0, 1'b1,  8'd11,    9'd0},
{  1'b0, 1'b0, 8'd156,    9'd0},{  1'b0, 1'b0, 8'd155,    9'd0},{  1'b0, 1'b0,  8'd81,   9'd77},{  1'b0, 1'b0,  8'd24,  9'd351},{  1'b0, 1'b0,  8'd15,   9'd52},{  1'b0, 1'b0,  8'd12,    9'd0},{  1'b0, 1'b1,   8'd7,  9'd253},
{  1'b0, 1'b0, 8'd157,    9'd0},{  1'b0, 1'b0, 8'd156,    9'd0},{  1'b0, 1'b0,  8'd49,   9'd30},{  1'b0, 1'b0,  8'd34,  9'd232},{  1'b0, 1'b0,  8'd30,  9'd271},{  1'b0, 1'b0,  8'd13,    9'd0},{  1'b0, 1'b1,   8'd9,  9'd246},
{  1'b0, 1'b0, 8'd158,    9'd0},{  1'b0, 1'b0, 8'd157,    9'd0},{  1'b0, 1'b0,  8'd43,   9'd58},{  1'b0, 1'b0,  8'd32,  9'd206},{  1'b0, 1'b0,  8'd31,  9'd247},{  1'b0, 1'b0,  8'd14,    9'd0},{  1'b0, 1'b1,   8'd6,  9'd195},
{  1'b0, 1'b0, 8'd159,    9'd0},{  1'b0, 1'b0, 8'd158,    9'd0},{  1'b0, 1'b0,  8'd84,   9'd88},{  1'b0, 1'b0,  8'd79,  9'd138},{  1'b0, 1'b0,  8'd26,  9'd126},{  1'b0, 1'b0,  8'd22,  9'd345},{  1'b0, 1'b1,  8'd15,    9'd0},
{  1'b0, 1'b0, 8'd160,    9'd0},{  1'b0, 1'b0, 8'd159,    9'd0},{  1'b0, 1'b0,  8'd32,  9'd137},{  1'b0, 1'b0,  8'd20,   9'd16},{  1'b0, 1'b0,  8'd16,    9'd0},{  1'b0, 1'b0,  8'd13,  9'd245},{  1'b0, 1'b1,   8'd1,  9'd264},
{  1'b0, 1'b0, 8'd161,    9'd0},{  1'b0, 1'b0, 8'd160,    9'd0},{  1'b0, 1'b0,  8'd28,   9'd62},{  1'b0, 1'b0,  8'd24,  9'd284},{  1'b0, 1'b0,  8'd17,    9'd0},{  1'b0, 1'b0,  8'd17,  9'd164},{  1'b0, 1'b1,   8'd2,  9'd274},
{  1'b0, 1'b0, 8'd162,    9'd0},{  1'b0, 1'b0, 8'd161,    9'd0},{  1'b0, 1'b0,  8'd53,  9'd224},{  1'b0, 1'b0,  8'd39,  9'd267},{  1'b0, 1'b0,  8'd34,  9'd173},{  1'b0, 1'b0,  8'd18,    9'd0},{  1'b0, 1'b1,   8'd2,    9'd8},
{  1'b0, 1'b0, 8'd163,    9'd0},{  1'b0, 1'b0, 8'd162,    9'd0},{  1'b0, 1'b0,  8'd62,  9'd216},{  1'b0, 1'b0,  8'd35,   9'd78},{  1'b0, 1'b0,  8'd27,  9'd330},{  1'b0, 1'b0,  8'd19,    9'd0},{  1'b0, 1'b1,  8'd18,  9'd184},
{  1'b0, 1'b0, 8'd164,    9'd0},{  1'b0, 1'b0, 8'd163,    9'd0},{  1'b0, 1'b0,  8'd75,  9'd130},{  1'b0, 1'b0,  8'd22,  9'd284},{  1'b0, 1'b0,  8'd20,    9'd0},{  1'b0, 1'b0,   8'd9,  9'd187},{  1'b0, 1'b1,   8'd9,  9'd305},
{  1'b0, 1'b0, 8'd165,    9'd0},{  1'b0, 1'b0, 8'd164,    9'd0},{  1'b0, 1'b0,  8'd77,   9'd14},{  1'b0, 1'b0,  8'd69,  9'd103},{  1'b0, 1'b0,  8'd23,  9'd352},{  1'b0, 1'b0,  8'd22,  9'd217},{  1'b0, 1'b1,  8'd21,    9'd0},
{  1'b0, 1'b0, 8'd166,    9'd0},{  1'b0, 1'b0, 8'd165,    9'd0},{  1'b0, 1'b0,  8'd54,  9'd273},{  1'b0, 1'b0,  8'd29,  9'd289},{  1'b0, 1'b0,  8'd26,  9'd242},{  1'b0, 1'b0,  8'd22,    9'd0},{  1'b0, 1'b1,  8'd14,  9'd203},
{  1'b0, 1'b0, 8'd167,    9'd0},{  1'b0, 1'b0, 8'd166,    9'd0},{  1'b0, 1'b0,  8'd36,  9'd161},{  1'b0, 1'b0,  8'd28,  9'd252},{  1'b0, 1'b0,  8'd24,  9'd256},{  1'b0, 1'b0,  8'd23,    9'd0},{  1'b0, 1'b1,   8'd7,  9'd125},
{  1'b0, 1'b0, 8'd168,    9'd0},{  1'b0, 1'b0, 8'd167,    9'd0},{  1'b0, 1'b0,  8'd44,  9'd312},{  1'b0, 1'b0,  8'd41,  9'd176},{  1'b0, 1'b0,  8'd24,    9'd0},{  1'b0, 1'b0,  8'd15,  9'd275},{  1'b0, 1'b1,  8'd13,  9'd151},
{  1'b0, 1'b0, 8'd169,    9'd0},{  1'b0, 1'b0, 8'd168,    9'd0},{  1'b0, 1'b0,  8'd82,   9'd10},{  1'b0, 1'b0,  8'd48,  9'd199},{  1'b0, 1'b0,  8'd25,    9'd0},{  1'b0, 1'b0,  8'd22,  9'd243},{  1'b0, 1'b1,   8'd2,  9'd101},
{  1'b0, 1'b0, 8'd170,    9'd0},{  1'b0, 1'b0, 8'd169,    9'd0},{  1'b0, 1'b0,  8'd80,  9'd356},{  1'b0, 1'b0,  8'd64,   9'd98},{  1'b0, 1'b0,  8'd26,    9'd0},{  1'b0, 1'b0,  8'd13,  9'd331},{  1'b0, 1'b1,   8'd2,   9'd63},
{  1'b0, 1'b0, 8'd171,    9'd0},{  1'b0, 1'b0, 8'd170,    9'd0},{  1'b0, 1'b0,  8'd76,  9'd333},{  1'b0, 1'b0,  8'd72,  9'd124},{  1'b0, 1'b0,  8'd34,  9'd253},{  1'b0, 1'b0,  8'd27,    9'd0},{  1'b0, 1'b1,  8'd16,  9'd243},
{  1'b0, 1'b0, 8'd172,    9'd0},{  1'b0, 1'b0, 8'd171,    9'd0},{  1'b0, 1'b0,  8'd55,  9'd354},{  1'b0, 1'b0,  8'd34,  9'd167},{  1'b0, 1'b0,  8'd28,    9'd0},{  1'b0, 1'b0,   8'd9,  9'd287},{  1'b0, 1'b1,   8'd0,  9'd159},
{  1'b0, 1'b0, 8'd173,    9'd0},{  1'b0, 1'b0, 8'd172,    9'd0},{  1'b0, 1'b0,  8'd62,   9'd15},{  1'b0, 1'b0,  8'd33,  9'd217},{  1'b0, 1'b0,  8'd29,    9'd0},{  1'b0, 1'b0,  8'd27,    9'd2},{  1'b0, 1'b1,   8'd7,  9'd157},
{  1'b0, 1'b0, 8'd174,    9'd0},{  1'b0, 1'b0, 8'd173,    9'd0},{  1'b0, 1'b0,  8'd69,  9'd329},{  1'b0, 1'b0,  8'd30,    9'd0},{  1'b0, 1'b0,  8'd28,  9'd242},{  1'b0, 1'b0,  8'd18,    9'd6},{  1'b0, 1'b1,  8'd11,  9'd189},
{  1'b0, 1'b0, 8'd175,    9'd0},{  1'b0, 1'b0, 8'd174,    9'd0},{  1'b0, 1'b0,  8'd33,   9'd66},{  1'b0, 1'b0,  8'd31,    9'd0},{  1'b0, 1'b0,  8'd29,  9'd334},{  1'b0, 1'b0,  8'd10,  9'd162},{  1'b0, 1'b1,   8'd9,  9'd237},
{  1'b0, 1'b0, 8'd176,    9'd0},{  1'b0, 1'b0, 8'd175,    9'd0},{  1'b0, 1'b0,  8'd32,    9'd0},{  1'b0, 1'b0,  8'd32,  9'd324},{  1'b0, 1'b0,  8'd31,  9'd336},{  1'b0, 1'b0,  8'd23,  9'd118},{  1'b0, 1'b1,   8'd8,  9'd332},
{  1'b0, 1'b0, 8'd177,    9'd0},{  1'b0, 1'b0, 8'd176,    9'd0},{  1'b0, 1'b0,  8'd84,  9'd241},{  1'b0, 1'b0,  8'd42,  9'd236},{  1'b0, 1'b0,  8'd33,    9'd0},{  1'b0, 1'b0,  8'd25,  9'd353},{  1'b0, 1'b1,  8'd11,  9'd259},
{  1'b0, 1'b0, 8'd178,    9'd0},{  1'b0, 1'b0, 8'd177,    9'd0},{  1'b0, 1'b0,  8'd56,  9'd221},{  1'b0, 1'b0,  8'd34,    9'd0},{  1'b0, 1'b0,  8'd15,  9'd153},{  1'b0, 1'b0,   8'd7,    9'd7},{  1'b0, 1'b1,   8'd5,  9'd177},
{  1'b0, 1'b0, 8'd179,    9'd0},{  1'b0, 1'b0, 8'd178,    9'd0},{  1'b0, 1'b0,  8'd43,  9'd161},{  1'b0, 1'b0,  8'd35,    9'd0},{  1'b0, 1'b0,  8'd32,  9'd358},{  1'b0, 1'b0,  8'd19,  9'd216},{  1'b0, 1'b1,   8'd0,  9'd298}
};
localparam bit [18 : 0] cLARGE_HS_V_TAB_1BY2_PACKED[cLARGE_HS_TAB_1BY2_PACKED_SIZE] = '{
{8'd179, 1'b0,   10'd0},{8'd179, 1'b1, 10'd623},
{8'd178, 1'b0, 10'd616},{8'd178, 1'b1, 10'd624},
{8'd177, 1'b0, 10'd609},{8'd177, 1'b1, 10'd617},
{8'd176, 1'b0, 10'd602},{8'd176, 1'b1, 10'd610},
{8'd175, 1'b0, 10'd595},{8'd175, 1'b1, 10'd603},
{8'd174, 1'b0, 10'd588},{8'd174, 1'b1, 10'd596},
{8'd173, 1'b0, 10'd581},{8'd173, 1'b1, 10'd589},
{8'd172, 1'b0, 10'd574},{8'd172, 1'b1, 10'd582},
{8'd171, 1'b0, 10'd567},{8'd171, 1'b1, 10'd575},
{8'd170, 1'b0, 10'd560},{8'd170, 1'b1, 10'd568},
{8'd169, 1'b0, 10'd553},{8'd169, 1'b1, 10'd561},
{8'd168, 1'b0, 10'd546},{8'd168, 1'b1, 10'd554},
{8'd167, 1'b0, 10'd539},{8'd167, 1'b1, 10'd547},
{8'd166, 1'b0, 10'd532},{8'd166, 1'b1, 10'd540},
{8'd165, 1'b0, 10'd525},{8'd165, 1'b1, 10'd533},
{8'd164, 1'b0, 10'd518},{8'd164, 1'b1, 10'd526},
{8'd163, 1'b0, 10'd511},{8'd163, 1'b1, 10'd519},
{8'd162, 1'b0, 10'd504},{8'd162, 1'b1, 10'd512},
{8'd161, 1'b0, 10'd497},{8'd161, 1'b1, 10'd505},
{8'd160, 1'b0, 10'd490},{8'd160, 1'b1, 10'd498},
{8'd159, 1'b0, 10'd483},{8'd159, 1'b1, 10'd491},
{8'd158, 1'b0, 10'd476},{8'd158, 1'b1, 10'd484},
{8'd157, 1'b0, 10'd469},{8'd157, 1'b1, 10'd477},
{8'd156, 1'b0, 10'd462},{8'd156, 1'b1, 10'd470},
{8'd155, 1'b0, 10'd455},{8'd155, 1'b1, 10'd463},
{8'd154, 1'b0, 10'd448},{8'd154, 1'b1, 10'd456},
{8'd153, 1'b0, 10'd441},{8'd153, 1'b1, 10'd449},
{8'd152, 1'b0, 10'd434},{8'd152, 1'b1, 10'd442},
{8'd151, 1'b0, 10'd427},{8'd151, 1'b1, 10'd435},
{8'd150, 1'b0, 10'd420},{8'd150, 1'b1, 10'd428},
{8'd149, 1'b0, 10'd413},{8'd149, 1'b1, 10'd421},
{8'd148, 1'b0, 10'd406},{8'd148, 1'b1, 10'd414},
{8'd147, 1'b0, 10'd399},{8'd147, 1'b1, 10'd407},
{8'd146, 1'b0, 10'd392},{8'd146, 1'b1, 10'd400},
{8'd145, 1'b0, 10'd385},{8'd145, 1'b1, 10'd393},
{8'd144, 1'b0, 10'd378},{8'd144, 1'b1, 10'd386},
{8'd143, 1'b0, 10'd371},{8'd143, 1'b1, 10'd379},
{8'd142, 1'b0, 10'd364},{8'd142, 1'b1, 10'd372},
{8'd141, 1'b0, 10'd357},{8'd141, 1'b1, 10'd365},
{8'd140, 1'b0, 10'd350},{8'd140, 1'b1, 10'd358},
{8'd139, 1'b0, 10'd343},{8'd139, 1'b1, 10'd351},
{8'd138, 1'b0, 10'd336},{8'd138, 1'b1, 10'd344},
{8'd137, 1'b0, 10'd329},{8'd137, 1'b1, 10'd337},
{8'd136, 1'b0, 10'd322},{8'd136, 1'b1, 10'd330},
{8'd135, 1'b0, 10'd315},{8'd135, 1'b1, 10'd323},
{8'd134, 1'b0, 10'd308},{8'd134, 1'b1, 10'd316},
{8'd133, 1'b0, 10'd301},{8'd133, 1'b1, 10'd309},
{8'd132, 1'b0, 10'd294},{8'd132, 1'b1, 10'd302},
{8'd131, 1'b0, 10'd287},{8'd131, 1'b1, 10'd295},
{8'd130, 1'b0, 10'd280},{8'd130, 1'b1, 10'd288},
{8'd129, 1'b0, 10'd273},{8'd129, 1'b1, 10'd281},
{8'd128, 1'b0, 10'd266},{8'd128, 1'b1, 10'd274},
{8'd127, 1'b0, 10'd259},{8'd127, 1'b1, 10'd267},
{8'd126, 1'b0, 10'd252},{8'd126, 1'b1, 10'd260},
{8'd125, 1'b0, 10'd245},{8'd125, 1'b1, 10'd253},
{8'd124, 1'b0, 10'd238},{8'd124, 1'b1, 10'd246},
{8'd123, 1'b0, 10'd231},{8'd123, 1'b1, 10'd239},
{8'd122, 1'b0, 10'd224},{8'd122, 1'b1, 10'd232},
{8'd121, 1'b0, 10'd217},{8'd121, 1'b1, 10'd225},
{8'd120, 1'b0, 10'd210},{8'd120, 1'b1, 10'd218},
{8'd119, 1'b0, 10'd203},{8'd119, 1'b1, 10'd211},
{8'd118, 1'b0, 10'd196},{8'd118, 1'b1, 10'd204},
{8'd117, 1'b0, 10'd189},{8'd117, 1'b1, 10'd197},
{8'd116, 1'b0, 10'd182},{8'd116, 1'b1, 10'd190},
{8'd115, 1'b0, 10'd175},{8'd115, 1'b1, 10'd183},
{8'd114, 1'b0, 10'd168},{8'd114, 1'b1, 10'd176},
{8'd113, 1'b0, 10'd161},{8'd113, 1'b1, 10'd169},
{8'd112, 1'b0, 10'd154},{8'd112, 1'b1, 10'd162},
{8'd111, 1'b0, 10'd147},{8'd111, 1'b1, 10'd155},
{8'd110, 1'b0, 10'd140},{8'd110, 1'b1, 10'd148},
{8'd109, 1'b0, 10'd133},{8'd109, 1'b1, 10'd141},
{8'd108, 1'b0, 10'd126},{8'd108, 1'b1, 10'd134},
{8'd107, 1'b0, 10'd119},{8'd107, 1'b1, 10'd127},
{8'd106, 1'b0, 10'd112},{8'd106, 1'b1, 10'd120},
{8'd105, 1'b0, 10'd105},{8'd105, 1'b1, 10'd113},
{8'd104, 1'b0,  10'd98},{8'd104, 1'b1, 10'd106},
{8'd103, 1'b0,  10'd91},{8'd103, 1'b1,  10'd99},
{8'd102, 1'b0,  10'd84},{8'd102, 1'b1,  10'd92},
{8'd101, 1'b0,  10'd77},{8'd101, 1'b1,  10'd85},
{8'd100, 1'b0,  10'd70},{8'd100, 1'b1,  10'd78},
{ 8'd99, 1'b0,  10'd63},{ 8'd99, 1'b1,  10'd71},
{ 8'd98, 1'b0,  10'd56},{ 8'd98, 1'b1,  10'd64},
{ 8'd97, 1'b0,  10'd49},{ 8'd97, 1'b1,  10'd57},
{ 8'd96, 1'b0,  10'd42},{ 8'd96, 1'b1,  10'd50},
{ 8'd95, 1'b0,  10'd35},{ 8'd95, 1'b1,  10'd43},
{ 8'd94, 1'b0,  10'd28},{ 8'd94, 1'b1,  10'd36},
{ 8'd93, 1'b0,  10'd21},{ 8'd93, 1'b1,  10'd29},
{ 8'd92, 1'b0,  10'd14},{ 8'd92, 1'b1,  10'd22},
{ 8'd91, 1'b0,   10'd7},{ 8'd91, 1'b1,  10'd15},
{ 8'd90, 1'b0,   10'd1},{ 8'd90, 1'b1,   10'd8},
{ 8'd89, 1'b0,  10'd51},{ 8'd89, 1'b0, 10'd303},{ 8'd89, 1'b1, 10'd373},
{ 8'd88, 1'b0, 10'd240},{ 8'd88, 1'b0, 10'd366},{ 8'd88, 1'b1, 10'd387},
{ 8'd87, 1'b0,  10'd58},{ 8'd87, 1'b0, 10'd359},{ 8'd87, 1'b1, 10'd367},
{ 8'd86, 1'b0, 10'd212},{ 8'd86, 1'b0, 10'd296},{ 8'd86, 1'b1, 10'd352},
{ 8'd85, 1'b0, 10'd156},{ 8'd85, 1'b0, 10'd345},{ 8'd85, 1'b1, 10'd360},
{ 8'd84, 1'b0, 10'd338},{ 8'd84, 1'b0, 10'd485},{ 8'd84, 1'b1, 10'd611},
{ 8'd83, 1'b0, 10'd184},{ 8'd83, 1'b0, 10'd331},{ 8'd83, 1'b1, 10'd380},
{ 8'd82, 1'b0,  10'd30},{ 8'd82, 1'b0, 10'd324},{ 8'd82, 1'b1, 10'd555},
{ 8'd81, 1'b0, 10'd128},{ 8'd81, 1'b0, 10'd317},{ 8'd81, 1'b1, 10'd464},
{ 8'd80, 1'b0, 10'd219},{ 8'd80, 1'b0, 10'd310},{ 8'd80, 1'b1, 10'd562},
{ 8'd79, 1'b0,  10'd65},{ 8'd79, 1'b0, 10'd304},{ 8'd79, 1'b1, 10'd486},
{ 8'd78, 1'b0,  10'd86},{ 8'd78, 1'b0, 10'd177},{ 8'd78, 1'b1, 10'd297},
{ 8'd77, 1'b0, 10'd241},{ 8'd77, 1'b0, 10'd289},{ 8'd77, 1'b1, 10'd527},
{ 8'd76, 1'b0,  10'd44},{ 8'd76, 1'b0, 10'd282},{ 8'd76, 1'b1, 10'd569},
{ 8'd75, 1'b0, 10'd275},{ 8'd75, 1'b0, 10'd283},{ 8'd75, 1'b1, 10'd520},
{ 8'd74, 1'b0,   10'd2},{ 8'd74, 1'b0, 10'd142},{ 8'd74, 1'b1, 10'd268},
{ 8'd73, 1'b0, 10'd114},{ 8'd73, 1'b0, 10'd261},{ 8'd73, 1'b1, 10'd368},
{ 8'd72, 1'b0, 10'd254},{ 8'd72, 1'b0, 10'd457},{ 8'd72, 1'b1, 10'd570},
{ 8'd71, 1'b0, 10'd157},{ 8'd71, 1'b0, 10'd247},{ 8'd71, 1'b1, 10'd325},
{ 8'd70, 1'b0, 10'd242},{ 8'd70, 1'b0, 10'd284},{ 8'd70, 1'b1, 10'd429},
{ 8'd69, 1'b0, 10'd233},{ 8'd69, 1'b0, 10'd528},{ 8'd69, 1'b1, 10'd590},
{ 8'd68, 1'b0,  10'd23},{ 8'd68, 1'b0, 10'd226},{ 8'd68, 1'b1, 10'd374},
{ 8'd67, 1'b0, 10'd100},{ 8'd67, 1'b0, 10'd149},{ 8'd67, 1'b1, 10'd220},
{ 8'd66, 1'b0,  10'd93},{ 8'd66, 1'b0, 10'd191},{ 8'd66, 1'b1, 10'd213},
{ 8'd65, 1'b0, 10'd205},{ 8'd65, 1'b0, 10'd332},{ 8'd65, 1'b1, 10'd436},
{ 8'd64, 1'b0, 10'd198},{ 8'd64, 1'b0, 10'd227},{ 8'd64, 1'b1, 10'd563},
{ 8'd63, 1'b0, 10'd101},{ 8'd63, 1'b0, 10'd107},{ 8'd63, 1'b1, 10'd192},
{ 8'd62, 1'b0, 10'd185},{ 8'd62, 1'b0, 10'd513},{ 8'd62, 1'b1, 10'd583},
{ 8'd61, 1'b0, 10'd178},{ 8'd61, 1'b0, 10'd262},{ 8'd61, 1'b1, 10'd430},
{ 8'd60, 1'b0, 10'd170},{ 8'd60, 1'b0, 10'd353},{ 8'd60, 1'b1, 10'd401},
{ 8'd59, 1'b0, 10'd115},{ 8'd59, 1'b0, 10'd163},{ 8'd59, 1'b1, 10'd305},
{ 8'd58, 1'b0,  10'd66},{ 8'd58, 1'b0, 10'd158},{ 8'd58, 1'b1, 10'd290},
{ 8'd57, 1'b0, 10'd150},{ 8'd57, 1'b0, 10'd291},{ 8'd57, 1'b1, 10'd422},
{ 8'd56, 1'b0, 10'd121},{ 8'd56, 1'b0, 10'd143},{ 8'd56, 1'b1, 10'd618},
{ 8'd55, 1'b0, 10'd135},{ 8'd55, 1'b0, 10'd276},{ 8'd55, 1'b1, 10'd576},
{ 8'd54, 1'b0, 10'd129},{ 8'd54, 1'b0, 10'd415},{ 8'd54, 1'b1, 10'd534},
{ 8'd53, 1'b0, 10'd122},{ 8'd53, 1'b0, 10'd388},{ 8'd53, 1'b1, 10'd506},
{ 8'd52, 1'b0, 10'd116},{ 8'd52, 1'b0, 10'd171},{ 8'd52, 1'b1, 10'd186},
{ 8'd51, 1'b0,  10'd16},{ 8'd51, 1'b0, 10'd108},{ 8'd51, 1'b1, 10'd255},
{ 8'd50, 1'b0, 10'd102},{ 8'd50, 1'b0, 10'd269},{ 8'd50, 1'b1, 10'd333},
{ 8'd49, 1'b0,  10'd94},{ 8'd49, 1'b0, 10'd123},{ 8'd49, 1'b1, 10'd471},
{ 8'd48, 1'b0,  10'd87},{ 8'd48, 1'b0, 10'd277},{ 8'd48, 1'b1, 10'd556},
{ 8'd47, 1'b0,  10'd79},{ 8'd47, 1'b0, 10'd214},{ 8'd47, 1'b1, 10'd458},
{ 8'd46, 1'b0,  10'd72},{ 8'd46, 1'b0,  10'd95},{ 8'd46, 1'b1, 10'd221},
{ 8'd45, 1'b0,  10'd67},{ 8'd45, 1'b0, 10'd164},{ 8'd45, 1'b1, 10'd199},
{ 8'd44, 1'b0,  10'd59},{ 8'd44, 1'b0, 10'd416},{ 8'd44, 1'b1, 10'd548},
{ 8'd43, 1'b0,  10'd52},{ 8'd43, 1'b0, 10'd478},{ 8'd43, 1'b1, 10'd625},
{ 8'd42, 1'b0,  10'd45},{ 8'd42, 1'b0, 10'd394},{ 8'd42, 1'b1, 10'd612},
{ 8'd41, 1'b0,   10'd9},{ 8'd41, 1'b0,  10'd37},{ 8'd41, 1'b1, 10'd549},
{ 8'd40, 1'b0,  10'd31},{ 8'd40, 1'b0, 10'd234},{ 8'd40, 1'b1, 10'd375},
{ 8'd39, 1'b0,  10'd24},{ 8'd39, 1'b0, 10'd311},{ 8'd39, 1'b1, 10'd507},
{ 8'd38, 1'b0,  10'd17},{ 8'd38, 1'b0, 10'd136},{ 8'd38, 1'b1, 10'd423},
{ 8'd37, 1'b0,  10'd10},{ 8'd37, 1'b0,  10'd73},{ 8'd37, 1'b1, 10'd270},
{ 8'd36, 1'b0,   10'd3},{ 8'd36, 1'b0, 10'd248},{ 8'd36, 1'b1, 10'd541},
{ 8'd35, 1'b0, 10'd172},{ 8'd35, 1'b0, 10'd206},{ 8'd35, 1'b0, 10'd235},{ 8'd35, 1'b0, 10'd339},{ 8'd35, 1'b0, 10'd408},{ 8'd35, 1'b0, 10'd437},{ 8'd35, 1'b0, 10'd514},{ 8'd35, 1'b1, 10'd626},
{ 8'd34, 1'b0,  10'd53},{ 8'd34, 1'b0, 10'd193},{ 8'd34, 1'b0, 10'd443},{ 8'd34, 1'b0, 10'd472},{ 8'd34, 1'b0, 10'd508},{ 8'd34, 1'b0, 10'd571},{ 8'd34, 1'b0, 10'd577},{ 8'd34, 1'b1, 10'd619},
{ 8'd33, 1'b0,  10'd32},{ 8'd33, 1'b0,  10'd88},{ 8'd33, 1'b0, 10'd326},{ 8'd33, 1'b0, 10'd346},{ 8'd33, 1'b0, 10'd450},{ 8'd33, 1'b0, 10'd584},{ 8'd33, 1'b0, 10'd597},{ 8'd33, 1'b1, 10'd613},
{ 8'd32, 1'b0,  10'd46},{ 8'd32, 1'b0,  10'd80},{ 8'd32, 1'b0, 10'd200},{ 8'd32, 1'b0, 10'd479},{ 8'd32, 1'b0, 10'd492},{ 8'd32, 1'b0, 10'd604},{ 8'd32, 1'b0, 10'd605},{ 8'd32, 1'b1, 10'd627},
{ 8'd31, 1'b0, 10'd144},{ 8'd31, 1'b0, 10'd159},{ 8'd31, 1'b0, 10'd263},{ 8'd31, 1'b0, 10'd292},{ 8'd31, 1'b0, 10'd431},{ 8'd31, 1'b0, 10'd480},{ 8'd31, 1'b0, 10'd598},{ 8'd31, 1'b1, 10'd606},
{ 8'd30, 1'b0,   10'd4},{ 8'd30, 1'b0,  10'd38},{ 8'd30, 1'b0,  10'd60},{ 8'd30, 1'b0, 10'd109},{ 8'd30, 1'b0, 10'd389},{ 8'd30, 1'b0, 10'd395},{ 8'd30, 1'b0, 10'd473},{ 8'd30, 1'b1, 10'd591},
{ 8'd29, 1'b0, 10'd187},{ 8'd29, 1'b0, 10'd347},{ 8'd29, 1'b0, 10'd409},{ 8'd29, 1'b0, 10'd417},{ 8'd29, 1'b0, 10'd444},{ 8'd29, 1'b0, 10'd535},{ 8'd29, 1'b0, 10'd585},{ 8'd29, 1'b1, 10'd599},
{ 8'd28, 1'b0,  10'd54},{ 8'd28, 1'b0, 10'd137},{ 8'd28, 1'b0, 10'd249},{ 8'd28, 1'b0, 10'd396},{ 8'd28, 1'b0, 10'd499},{ 8'd28, 1'b0, 10'd542},{ 8'd28, 1'b0, 10'd578},{ 8'd28, 1'b1, 10'd592},
{ 8'd27, 1'b0,   10'd5},{ 8'd27, 1'b0,  10'd18},{ 8'd27, 1'b0, 10'd124},{ 8'd27, 1'b0, 10'd179},{ 8'd27, 1'b0, 10'd298},{ 8'd27, 1'b0, 10'd515},{ 8'd27, 1'b0, 10'd572},{ 8'd27, 1'b1, 10'd586},
{ 8'd26, 1'b0,   10'd6},{ 8'd26, 1'b0,  10'd89},{ 8'd26, 1'b0, 10'd278},{ 8'd26, 1'b0, 10'd334},{ 8'd26, 1'b0, 10'd402},{ 8'd26, 1'b0, 10'd487},{ 8'd26, 1'b0, 10'd536},{ 8'd26, 1'b1, 10'd564},
{ 8'd25, 1'b0, 10'd130},{ 8'd25, 1'b0, 10'd201},{ 8'd25, 1'b0, 10'd228},{ 8'd25, 1'b0, 10'd256},{ 8'd25, 1'b0, 10'd312},{ 8'd25, 1'b0, 10'd390},{ 8'd25, 1'b0, 10'd557},{ 8'd25, 1'b1, 10'd614},
{ 8'd24, 1'b0,  10'd33},{ 8'd24, 1'b0,  10'd39},{ 8'd24, 1'b0,  10'd68},{ 8'd24, 1'b0, 10'd180},{ 8'd24, 1'b0, 10'd465},{ 8'd24, 1'b0, 10'd500},{ 8'd24, 1'b0, 10'd543},{ 8'd24, 1'b1, 10'd550},
{ 8'd23, 1'b0, 10'd110},{ 8'd23, 1'b0, 10'd131},{ 8'd23, 1'b0, 10'd376},{ 8'd23, 1'b0, 10'd410},{ 8'd23, 1'b0, 10'd451},{ 8'd23, 1'b0, 10'd529},{ 8'd23, 1'b0, 10'd544},{ 8'd23, 1'b1, 10'd607},
{ 8'd22, 1'b0, 10'd215},{ 8'd22, 1'b0, 10'd250},{ 8'd22, 1'b0, 10'd318},{ 8'd22, 1'b0, 10'd488},{ 8'd22, 1'b0, 10'd521},{ 8'd22, 1'b0, 10'd530},{ 8'd22, 1'b0, 10'd537},{ 8'd22, 1'b1, 10'd558},
{ 8'd21, 1'b0,  10'd47},{ 8'd21, 1'b0,  10'd69},{ 8'd21, 1'b0, 10'd257},{ 8'd21, 1'b0, 10'd306},{ 8'd21, 1'b0, 10'd327},{ 8'd21, 1'b0, 10'd361},{ 8'd21, 1'b0, 10'd424},{ 8'd21, 1'b1, 10'd531},
{ 8'd20, 1'b0,  10'd11},{ 8'd20, 1'b0,  10'd81},{ 8'd20, 1'b0, 10'd216},{ 8'd20, 1'b0, 10'd279},{ 8'd20, 1'b0, 10'd285},{ 8'd20, 1'b0, 10'd299},{ 8'd20, 1'b0, 10'd493},{ 8'd20, 1'b1, 10'd522},
{ 8'd19, 1'b0,  10'd82},{ 8'd19, 1'b0, 10'd145},{ 8'd19, 1'b0, 10'd160},{ 8'd19, 1'b0, 10'd165},{ 8'd19, 1'b0, 10'd181},{ 8'd19, 1'b0, 10'd313},{ 8'd19, 1'b0, 10'd516},{ 8'd19, 1'b1, 10'd628},
{ 8'd18, 1'b0,  10'd61},{ 8'd18, 1'b0, 10'd103},{ 8'd18, 1'b0, 10'd202},{ 8'd18, 1'b0, 10'd319},{ 8'd18, 1'b0, 10'd452},{ 8'd18, 1'b0, 10'd509},{ 8'd18, 1'b0, 10'd517},{ 8'd18, 1'b1, 10'd593},
{ 8'd17, 1'b0, 10'd173},{ 8'd17, 1'b0, 10'd229},{ 8'd17, 1'b0, 10'd293},{ 8'd17, 1'b0, 10'd369},{ 8'd17, 1'b0, 10'd418},{ 8'd17, 1'b0, 10'd459},{ 8'd17, 1'b0, 10'd501},{ 8'd17, 1'b1, 10'd502},
{ 8'd16, 1'b0,  10'd19},{ 8'd16, 1'b0,  10'd25},{ 8'd16, 1'b0,  10'd62},{ 8'd16, 1'b0,  10'd96},{ 8'd16, 1'b0, 10'd236},{ 8'd16, 1'b0, 10'd300},{ 8'd16, 1'b0, 10'd494},{ 8'd16, 1'b1, 10'd573},
{ 8'd15, 1'b0,  10'd90},{ 8'd15, 1'b0, 10'd138},{ 8'd15, 1'b0, 10'd237},{ 8'd15, 1'b0, 10'd286},{ 8'd15, 1'b0, 10'd466},{ 8'd15, 1'b0, 10'd489},{ 8'd15, 1'b0, 10'd551},{ 8'd15, 1'b1, 10'd620},
{ 8'd14, 1'b0,  10'd48},{ 8'd14, 1'b0, 10'd132},{ 8'd14, 1'b0, 10'd207},{ 8'd14, 1'b0, 10'd251},{ 8'd14, 1'b0, 10'd307},{ 8'd14, 1'b0, 10'd340},{ 8'd14, 1'b0, 10'd481},{ 8'd14, 1'b1, 10'd538},
{ 8'd13, 1'b0,  10'd40},{ 8'd13, 1'b0, 10'd111},{ 8'd13, 1'b0, 10'd194},{ 8'd13, 1'b0, 10'd460},{ 8'd13, 1'b0, 10'd474},{ 8'd13, 1'b0, 10'd495},{ 8'd13, 1'b0, 10'd552},{ 8'd13, 1'b1, 10'd565},
{ 8'd12, 1'b0, 10'd243},{ 8'd12, 1'b0, 10'd354},{ 8'd12, 1'b0, 10'd403},{ 8'd12, 1'b0, 10'd425},{ 8'd12, 1'b0, 10'd432},{ 8'd12, 1'b0, 10'd438},{ 8'd12, 1'b0, 10'd439},{ 8'd12, 1'b1, 10'd467},
{ 8'd11, 1'b0, 10'd117},{ 8'd11, 1'b0, 10'd146},{ 8'd11, 1'b0, 10'd151},{ 8'd11, 1'b0, 10'd244},{ 8'd11, 1'b0, 10'd355},{ 8'd11, 1'b0, 10'd461},{ 8'd11, 1'b0, 10'd594},{ 8'd11, 1'b1, 10'd615},
{ 8'd10, 1'b0,  10'd12},{ 8'd10, 1'b0,  10'd13},{ 8'd10, 1'b0, 10'd264},{ 8'd10, 1'b0, 10'd271},{ 8'd10, 1'b0, 10'd341},{ 8'd10, 1'b0, 10'd377},{ 8'd10, 1'b0, 10'd453},{ 8'd10, 1'b1, 10'd600},
{  8'd9, 1'b0,  10'd34},{  8'd9, 1'b0, 10'd166},{  8'd9, 1'b0, 10'd445},{  8'd9, 1'b0, 10'd475},{  8'd9, 1'b0, 10'd523},{  8'd9, 1'b0, 10'd524},{  8'd9, 1'b0, 10'd579},{  8'd9, 1'b1, 10'd601},
{  8'd8, 1'b0,  10'd83},{  8'd8, 1'b0,  10'd97},{  8'd8, 1'b0, 10'd125},{  8'd8, 1'b0, 10'd152},{  8'd8, 1'b0, 10'd314},{  8'd8, 1'b0, 10'd381},{  8'd8, 1'b0, 10'd440},{  8'd8, 1'b1, 10'd608},
{  8'd7, 1'b0, 10'd195},{  8'd7, 1'b0, 10'd272},{  8'd7, 1'b0, 10'd328},{  8'd7, 1'b0, 10'd433},{  8'd7, 1'b0, 10'd468},{  8'd7, 1'b0, 10'd545},{  8'd7, 1'b0, 10'd587},{  8'd7, 1'b1, 10'd621},
{  8'd6, 1'b0,  10'd26},{  8'd6, 1'b0, 10'd118},{  8'd6, 1'b0, 10'd208},{  8'd6, 1'b0, 10'd230},{  8'd6, 1'b0, 10'd382},{  8'd6, 1'b0, 10'd397},{  8'd6, 1'b0, 10'd426},{  8'd6, 1'b1, 10'd482},
{  8'd5, 1'b0,  10'd74},{  8'd5, 1'b0, 10'd209},{  8'd5, 1'b0, 10'd258},{  8'd5, 1'b0, 10'd320},{  8'd5, 1'b0, 10'd348},{  8'd5, 1'b0, 10'd370},{  8'd5, 1'b0, 10'd419},{  8'd5, 1'b1, 10'd622},
{  8'd4, 1'b0,  10'd20},{  8'd4, 1'b0,  10'd55},{  8'd4, 1'b0,  10'd75},{  8'd4, 1'b0, 10'd174},{  8'd4, 1'b0, 10'd222},{  8'd4, 1'b0, 10'd265},{  8'd4, 1'b0, 10'd411},{  8'd4, 1'b1, 10'd412},
{  8'd3, 1'b0,  10'd41},{  8'd3, 1'b0, 10'd167},{  8'd3, 1'b0, 10'd223},{  8'd3, 1'b0, 10'd362},{  8'd3, 1'b0, 10'd383},{  8'd3, 1'b0, 10'd404},{  8'd3, 1'b0, 10'd405},{  8'd3, 1'b1, 10'd454},
{  8'd2, 1'b0,  10'd27},{  8'd2, 1'b0, 10'd139},{  8'd2, 1'b0, 10'd188},{  8'd2, 1'b0, 10'd398},{  8'd2, 1'b0, 10'd503},{  8'd2, 1'b0, 10'd510},{  8'd2, 1'b0, 10'd559},{  8'd2, 1'b1, 10'd566},
{  8'd1, 1'b0,  10'd76},{  8'd1, 1'b0, 10'd321},{  8'd1, 1'b0, 10'd356},{  8'd1, 1'b0, 10'd363},{  8'd1, 1'b0, 10'd391},{  8'd1, 1'b0, 10'd446},{  8'd1, 1'b0, 10'd447},{  8'd1, 1'b1, 10'd496},
{  8'd0, 1'b0, 10'd104},{  8'd0, 1'b0, 10'd153},{  8'd0, 1'b0, 10'd335},{  8'd0, 1'b0, 10'd342},{  8'd0, 1'b0, 10'd349},{  8'd0, 1'b0, 10'd384},{  8'd0, 1'b0, 10'd580},{  8'd0, 1'b1, 10'd629}
};
localparam int          cLARGE_HS_TAB_3BY5_PACKED_SIZE = 792;
localparam bit [18 : 0] cLARGE_HS_TAB_3BY5_PACKED[cLARGE_HS_TAB_3BY5_PACKED_SIZE] = '{
{  1'b1, 1'b0, 8'd179,    9'd1},{  1'b0, 1'b0, 8'd108,    9'd0},{  1'b0, 1'b0, 8'd101,  9'd203},{  1'b0, 1'b0,  8'd40,  9'd209},{  1'b0, 1'b0,  8'd36,    9'd0},{  1'b0, 1'b0,  8'd33,  9'd114},{  1'b0, 1'b0,  8'd32,  9'd345},{  1'b0, 1'b0,  8'd24,  9'd134},{  1'b0, 1'b0,  8'd22,  9'd313},{  1'b0, 1'b0,  8'd15,  9'd200},{  1'b0, 1'b1,   8'd0,  9'd237},
{  1'b0, 1'b0, 8'd109,    9'd0},{  1'b0, 1'b0, 8'd108,    9'd0},{  1'b0, 1'b0,  8'd97,  9'd346},{  1'b0, 1'b0,  8'd44,   9'd74},{  1'b0, 1'b0,  8'd37,    9'd0},{  1'b0, 1'b0,  8'd33,  9'd134},{  1'b0, 1'b0,  8'd24,   9'd67},{  1'b0, 1'b0,  8'd11,  9'd262},{  1'b0, 1'b0,   8'd9,   9'd26},{  1'b0, 1'b0,   8'd7,  9'd138},{  1'b0, 1'b1,   8'd0,  9'd155},
{  1'b0, 1'b0, 8'd110,    9'd0},{  1'b0, 1'b0, 8'd109,    9'd0},{  1'b0, 1'b0,  8'd92,  9'd339},{  1'b0, 1'b0,  8'd64,   9'd94},{  1'b0, 1'b0,  8'd38,    9'd0},{  1'b0, 1'b0,  8'd34,   9'd35},{  1'b0, 1'b0,  8'd33,  9'd156},{  1'b0, 1'b0,  8'd14,   9'd52},{  1'b0, 1'b0,   8'd8,  9'd178},{  1'b0, 1'b0,   8'd6,  9'd257},{  1'b0, 1'b1,   8'd2,  9'd357},
{  1'b0, 1'b0, 8'd111,    9'd0},{  1'b0, 1'b0, 8'd110,    9'd0},{  1'b0, 1'b0, 8'd104,  9'd211},{  1'b0, 1'b0,  8'd57,  9'd359},{  1'b0, 1'b0,  8'd39,    9'd0},{  1'b0, 1'b0,  8'd27,  9'd243},{  1'b0, 1'b0,  8'd26,  9'd259},{  1'b0, 1'b0,  8'd22,  9'd145},{  1'b0, 1'b0,  8'd17,  9'd217},{  1'b0, 1'b0,  8'd17,  9'd186},{  1'b0, 1'b1,  8'd12,  9'd327},
{  1'b0, 1'b0, 8'd112,    9'd0},{  1'b0, 1'b0, 8'd111,    9'd0},{  1'b0, 1'b0,  8'd96,  9'd358},{  1'b0, 1'b0,  8'd55,   9'd23},{  1'b0, 1'b0,  8'd40,    9'd0},{  1'b0, 1'b0,  8'd25,   9'd34},{  1'b0, 1'b0,  8'd18,   9'd50},{  1'b0, 1'b0,  8'd18,  9'd121},{  1'b0, 1'b0,  8'd14,  9'd139},{  1'b0, 1'b0,  8'd11,  9'd125},{  1'b0, 1'b1,   8'd7,  9'd353},
{  1'b0, 1'b0, 8'd113,    9'd0},{  1'b0, 1'b0, 8'd112,    9'd0},{  1'b0, 1'b0,  8'd94,  9'd137},{  1'b0, 1'b0,  8'd48,  9'd201},{  1'b0, 1'b0,  8'd41,    9'd0},{  1'b0, 1'b0,  8'd31,  9'd120},{  1'b0, 1'b0,  8'd29,   9'd53},{  1'b0, 1'b0,  8'd28,   9'd11},{  1'b0, 1'b0,  8'd25,  9'd160},{  1'b0, 1'b0,  8'd24,  9'd210},{  1'b0, 1'b1,  8'd22,  9'd209},
{  1'b0, 1'b0, 8'd114,    9'd0},{  1'b0, 1'b0, 8'd113,    9'd0},{  1'b0, 1'b0,  8'd98,  9'd341},{  1'b0, 1'b0,  8'd50,  9'd184},{  1'b0, 1'b0,  8'd42,    9'd0},{  1'b0, 1'b0,  8'd25,  9'd285},{  1'b0, 1'b0,  8'd20,  9'd245},{  1'b0, 1'b0,  8'd17,  9'd352},{  1'b0, 1'b0,  8'd12,  9'd100},{  1'b0, 1'b0,  8'd10,  9'd180},{  1'b0, 1'b1,   8'd6,   9'd85},
{  1'b0, 1'b0, 8'd115,    9'd0},{  1'b0, 1'b0, 8'd114,    9'd0},{  1'b0, 1'b0,  8'd97,  9'd287},{  1'b0, 1'b0,  8'd45,  9'd259},{  1'b0, 1'b0,  8'd43,    9'd0},{  1'b0, 1'b0,  8'd31,   9'd44},{  1'b0, 1'b0,  8'd30,   9'd86},{  1'b0, 1'b0,  8'd27,  9'd298},{  1'b0, 1'b0,  8'd25,  9'd184},{  1'b0, 1'b0,  8'd18,  9'd228},{  1'b0, 1'b1,  8'd10,   9'd62},
{  1'b0, 1'b0, 8'd116,    9'd0},{  1'b0, 1'b0, 8'd115,    9'd0},{  1'b0, 1'b0,  8'd79,  9'd357},{  1'b0, 1'b0,  8'd44,    9'd0},{  1'b0, 1'b0,  8'd38,  9'd130},{  1'b0, 1'b0,  8'd35,  9'd246},{  1'b0, 1'b0,  8'd22,   9'd56},{  1'b0, 1'b0,   8'd8,   9'd88},{  1'b0, 1'b0,   8'd8,   9'd98},{  1'b0, 1'b0,   8'd8,  9'd121},{  1'b0, 1'b1,   8'd3,  9'd354},
{  1'b0, 1'b0, 8'd117,    9'd0},{  1'b0, 1'b0, 8'd116,    9'd0},{  1'b0, 1'b0,  8'd77,  9'd342},{  1'b0, 1'b0,  8'd67,   9'd64},{  1'b0, 1'b0,  8'd45,    9'd0},{  1'b0, 1'b0,  8'd31,  9'd169},{  1'b0, 1'b0,  8'd30,  9'd329},{  1'b0, 1'b0,  8'd22,   9'd66},{  1'b0, 1'b0,  8'd11,  9'd157},{  1'b0, 1'b0,   8'd7,  9'd117},{  1'b0, 1'b1,   8'd0,   9'd78},
{  1'b0, 1'b0, 8'd118,    9'd0},{  1'b0, 1'b0, 8'd117,    9'd0},{  1'b0, 1'b0, 8'd103,   9'd13},{  1'b0, 1'b0,  8'd51,  9'd267},{  1'b0, 1'b0,  8'd46,    9'd0},{  1'b0, 1'b0,  8'd30,  9'd131},{  1'b0, 1'b0,  8'd24,  9'd234},{  1'b0, 1'b0,  8'd23,  9'd187},{  1'b0, 1'b0,  8'd17,   9'd81},{  1'b0, 1'b0,  8'd13,   9'd61},{  1'b0, 1'b1,   8'd1,   9'd58},
{  1'b0, 1'b0, 8'd119,    9'd0},{  1'b0, 1'b0, 8'd118,    9'd0},{  1'b0, 1'b0,  8'd82,  9'd288},{  1'b0, 1'b0,  8'd56,   9'd61},{  1'b0, 1'b0,  8'd47,    9'd0},{  1'b0, 1'b0,  8'd16,  9'd243},{  1'b0, 1'b0,  8'd15,  9'd336},{  1'b0, 1'b0,  8'd11,   9'd92},{  1'b0, 1'b0,  8'd11,  9'd136},{  1'b0, 1'b0,   8'd9,  9'd300},{  1'b0, 1'b1,   8'd4,  9'd106},
{  1'b0, 1'b0, 8'd120,    9'd0},{  1'b0, 1'b0, 8'd119,    9'd0},{  1'b0, 1'b0,  8'd94,  9'd114},{  1'b0, 1'b0,  8'd48,    9'd0},{  1'b0, 1'b0,  8'd41,  9'd256},{  1'b0, 1'b0,  8'd35,  9'd103},{  1'b0, 1'b0,  8'd33,  9'd346},{  1'b0, 1'b0,  8'd25,  9'd280},{  1'b0, 1'b0,  8'd13,  9'd162},{  1'b0, 1'b0,  8'd11,  9'd202},{  1'b0, 1'b1,   8'd5,   9'd74},
{  1'b0, 1'b0, 8'd121,    9'd0},{  1'b0, 1'b0, 8'd120,    9'd0},{  1'b0, 1'b0,  8'd81,   9'd14},{  1'b0, 1'b0,  8'd49,    9'd0},{  1'b0, 1'b0,  8'd36,  9'd259},{  1'b0, 1'b0,  8'd34,  9'd163},{  1'b0, 1'b0,  8'd31,   9'd40},{  1'b0, 1'b0,  8'd15,  9'd319},{  1'b0, 1'b0,   8'd7,   9'd51},{  1'b0, 1'b0,   8'd3,   9'd95},{  1'b0, 1'b1,   8'd3,  9'd221},
{  1'b0, 1'b0, 8'd122,    9'd0},{  1'b0, 1'b0, 8'd121,    9'd0},{  1'b0, 1'b0,  8'd89,   9'd96},{  1'b0, 1'b0,  8'd69,   9'd28},{  1'b0, 1'b0,  8'd50,    9'd0},{  1'b0, 1'b0,  8'd29,  9'd352},{  1'b0, 1'b0,  8'd28,  9'd318},{  1'b0, 1'b0,  8'd17,  9'd332},{  1'b0, 1'b0,  8'd15,  9'd111},{  1'b0, 1'b0,  8'd13,  9'd285},{  1'b0, 1'b1,   8'd7,   9'd65},
{  1'b0, 1'b0, 8'd123,    9'd0},{  1'b0, 1'b0, 8'd122,    9'd0},{  1'b0, 1'b0,  8'd80,  9'd167},{  1'b0, 1'b0,  8'd60,  9'd223},{  1'b0, 1'b0,  8'd51,    9'd0},{  1'b0, 1'b0,  8'd32,  9'd117},{  1'b0, 1'b0,  8'd31,  9'd143},{  1'b0, 1'b0,  8'd27,  9'd226},{  1'b0, 1'b0,  8'd23,  9'd306},{  1'b0, 1'b0,  8'd15,  9'd105},{  1'b0, 1'b1,   8'd4,  9'd201},
{  1'b0, 1'b0, 8'd124,    9'd0},{  1'b0, 1'b0, 8'd123,    9'd0},{  1'b0, 1'b0, 8'd102,   9'd51},{  1'b0, 1'b0,  8'd52,    9'd0},{  1'b0, 1'b0,  8'd41,  9'd342},{  1'b0, 1'b0,  8'd29,   9'd70},{  1'b0, 1'b0,  8'd27,  9'd262},{  1'b0, 1'b0,  8'd19,  9'd256},{  1'b0, 1'b0,  8'd15,   9'd71},{  1'b0, 1'b0,  8'd13,  9'd246},{  1'b0, 1'b1,   8'd9,  9'd321},
{  1'b0, 1'b0, 8'd125,    9'd0},{  1'b0, 1'b0, 8'd124,    9'd0},{  1'b0, 1'b0,  8'd90,   9'd86},{  1'b0, 1'b0,  8'd60,  9'd300},{  1'b0, 1'b0,  8'd53,    9'd0},{  1'b0, 1'b0,  8'd35,   9'd88},{  1'b0, 1'b0,  8'd29,  9'd319},{  1'b0, 1'b0,  8'd26,  9'd204},{  1'b0, 1'b0,  8'd23,    9'd5},{  1'b0, 1'b0,   8'd5,  9'd352},{  1'b0, 1'b1,   8'd2,   9'd30},
{  1'b0, 1'b0, 8'd126,    9'd0},{  1'b0, 1'b0, 8'd125,    9'd0},{  1'b0, 1'b0,  8'd99,  9'd172},{  1'b0, 1'b0,  8'd58,  9'd316},{  1'b0, 1'b0,  8'd54,    9'd0},{  1'b0, 1'b0,  8'd23,  9'd336},{  1'b0, 1'b0,  8'd20,   9'd84},{  1'b0, 1'b0,  8'd14,  9'd129},{  1'b0, 1'b0,  8'd14,   9'd40},{  1'b0, 1'b0,   8'd4,  9'd242},{  1'b0, 1'b1,   8'd1,  9'd225},
{  1'b0, 1'b0, 8'd127,    9'd0},{  1'b0, 1'b0, 8'd126,    9'd0},{  1'b0, 1'b0,  8'd91,  9'd193},{  1'b0, 1'b0,  8'd59,  9'd196},{  1'b0, 1'b0,  8'd55,    9'd0},{  1'b0, 1'b0,  8'd31,   9'd51},{  1'b0, 1'b0,  8'd27,   9'd41},{  1'b0, 1'b0,   8'd9,  9'd104},{  1'b0, 1'b0,   8'd7,  9'd356},{  1'b0, 1'b0,   8'd5,   9'd78},{  1'b0, 1'b1,   8'd2,  9'd188},
{  1'b0, 1'b0, 8'd128,    9'd0},{  1'b0, 1'b0, 8'd127,    9'd0},{  1'b0, 1'b0,  8'd92,  9'd183},{  1'b0, 1'b0,  8'd63,  9'd112},{  1'b0, 1'b0,  8'd56,    9'd0},{  1'b0, 1'b0,  8'd32,  9'd304},{  1'b0, 1'b0,  8'd23,  9'd166},{  1'b0, 1'b0,  8'd19,  9'd122},{  1'b0, 1'b0,  8'd11,  9'd307},{  1'b0, 1'b0,  8'd10,  9'd290},{  1'b0, 1'b1,   8'd2,  9'd121},
{  1'b0, 1'b0, 8'd129,    9'd0},{  1'b0, 1'b0, 8'd128,    9'd0},{  1'b0, 1'b0,  8'd75,   9'd71},{  1'b0, 1'b0,  8'd62,    9'd8},{  1'b0, 1'b0,  8'd57,    9'd0},{  1'b0, 1'b0,  8'd18,  9'd227},{  1'b0, 1'b0,  8'd15,  9'd181},{  1'b0, 1'b0,   8'd6,   9'd75},{  1'b0, 1'b0,   8'd4,  9'd336},{  1'b0, 1'b0,   8'd3,  9'd230},{  1'b0, 1'b1,   8'd2,  9'd267},
{  1'b0, 1'b0, 8'd130,    9'd0},{  1'b0, 1'b0, 8'd129,    9'd0},{  1'b0, 1'b0, 8'd102,  9'd236},{  1'b0, 1'b0,  8'd58,    9'd0},{  1'b0, 1'b0,  8'd49,   9'd10},{  1'b0, 1'b0,  8'd29,  9'd264},{  1'b0, 1'b0,  8'd26,  9'd211},{  1'b0, 1'b0,  8'd26,  9'd141},{  1'b0, 1'b0,  8'd21,  9'd230},{  1'b0, 1'b0,  8'd17,   9'd58},{  1'b0, 1'b1,   8'd3,  9'd302},
{  1'b0, 1'b0, 8'd131,    9'd0},{  1'b0, 1'b0, 8'd130,    9'd0},{  1'b0, 1'b0,  8'd79,  9'd304},{  1'b0, 1'b0,  8'd59,    9'd0},{  1'b0, 1'b0,  8'd42,  9'd266},{  1'b0, 1'b0,  8'd27,   9'd57},{  1'b0, 1'b0,  8'd27,  9'd110},{  1'b0, 1'b0,  8'd27,   9'd77},{  1'b0, 1'b0,  8'd19,  9'd289},{  1'b0, 1'b0,   8'd9,  9'd285},{  1'b0, 1'b1,   8'd1,  9'd236},
{  1'b0, 1'b0, 8'd132,    9'd0},{  1'b0, 1'b0, 8'd131,    9'd0},{  1'b0, 1'b0,  8'd86,   9'd90},{  1'b0, 1'b0,  8'd62,  9'd277},{  1'b0, 1'b0,  8'd60,    9'd0},{  1'b0, 1'b0,  8'd35,   9'd34},{  1'b0, 1'b0,  8'd30,  9'd306},{  1'b0, 1'b0,  8'd21,  9'd338},{  1'b0, 1'b0,  8'd20,   9'd62},{  1'b0, 1'b0,   8'd6,  9'd124},{  1'b0, 1'b1,   8'd1,  9'd356},
{  1'b0, 1'b0, 8'd133,    9'd0},{  1'b0, 1'b0, 8'd132,    9'd0},{  1'b0, 1'b0,  8'd76,  9'd315},{  1'b0, 1'b0,  8'd61,    9'd0},{  1'b0, 1'b0,  8'd51,  9'd184},{  1'b0, 1'b0,  8'd32,  9'd284},{  1'b0, 1'b0,  8'd25,   9'd49},{  1'b0, 1'b0,  8'd17,  9'd207},{  1'b0, 1'b0,  8'd11,  9'd176},{  1'b0, 1'b0,   8'd1,  9'd278},{  1'b0, 1'b1,   8'd1,  9'd240},
{  1'b0, 1'b0, 8'd134,    9'd0},{  1'b0, 1'b0, 8'd133,    9'd0},{  1'b0, 1'b0,  8'd76,   9'd96},{  1'b0, 1'b0,  8'd62,    9'd0},{  1'b0, 1'b0,  8'd52,  9'd293},{  1'b0, 1'b0,  8'd35,   9'd21},{  1'b0, 1'b0,  8'd28,  9'd284},{  1'b0, 1'b0,  8'd17,  9'd212},{  1'b0, 1'b0,  8'd16,   9'd48},{  1'b0, 1'b0,  8'd14,  9'd275},{  1'b0, 1'b1,   8'd0,   9'd43},
{  1'b0, 1'b0, 8'd135,    9'd0},{  1'b0, 1'b0, 8'd134,    9'd0},{  1'b0, 1'b0,  8'd83,  9'd211},{  1'b0, 1'b0,  8'd63,    9'd0},{  1'b0, 1'b0,  8'd43,  9'd152},{  1'b0, 1'b0,  8'd35,   9'd50},{  1'b0, 1'b0,  8'd32,   9'd51},{  1'b0, 1'b0,  8'd16,  9'd181},{  1'b0, 1'b0,  8'd10,  9'd207},{  1'b0, 1'b0,   8'd6,  9'd181},{  1'b0, 1'b1,   8'd0,    9'd1},
{  1'b0, 1'b0, 8'd136,    9'd0},{  1'b0, 1'b0, 8'd135,    9'd0},{  1'b0, 1'b0,  8'd72,  9'd347},{  1'b0, 1'b0,  8'd64,    9'd0},{  1'b0, 1'b0,  8'd47,  9'd101},{  1'b0, 1'b0,  8'd32,  9'd253},{  1'b0, 1'b0,  8'd30,  9'd314},{  1'b0, 1'b0,  8'd18,  9'd133},{  1'b0, 1'b0,  8'd10,   9'd64},{  1'b0, 1'b0,  8'd10,  9'd171},{  1'b0, 1'b1,   8'd2,   9'd76},
{  1'b0, 1'b0, 8'd137,    9'd0},{  1'b0, 1'b0, 8'd136,    9'd0},{  1'b0, 1'b0,  8'd75,  9'd294},{  1'b0, 1'b0,  8'd65,    9'd0},{  1'b0, 1'b0,  8'd59,  9'd149},{  1'b0, 1'b0,  8'd30,  9'd228},{  1'b0, 1'b0,  8'd27,   9'd94},{  1'b0, 1'b0,  8'd11,  9'd311},{  1'b0, 1'b0,  8'd10,  9'd228},{  1'b0, 1'b0,   8'd5,  9'd280},{  1'b0, 1'b1,   8'd2,  9'd317},
{  1'b0, 1'b0, 8'd138,    9'd0},{  1'b0, 1'b0, 8'd137,    9'd0},{  1'b0, 1'b0,  8'd99,   9'd51},{  1'b0, 1'b0,  8'd66,    9'd0},{  1'b0, 1'b0,  8'd53,  9'd316},{  1'b0, 1'b0,  8'd29,  9'd329},{  1'b0, 1'b0,  8'd22,  9'd353},{  1'b0, 1'b0,  8'd13,  9'd203},{  1'b0, 1'b0,   8'd8,  9'd241},{  1'b0, 1'b0,   8'd8,   9'd73},{  1'b0, 1'b1,   8'd0,  9'd311},
{  1'b0, 1'b0, 8'd139,    9'd0},{  1'b0, 1'b0, 8'd138,    9'd0},{  1'b0, 1'b0,  8'd85,  9'd199},{  1'b0, 1'b0,  8'd67,    9'd0},{  1'b0, 1'b0,  8'd52,   9'd84},{  1'b0, 1'b0,  8'd33,  9'd150},{  1'b0, 1'b0,  8'd32,   9'd75},{  1'b0, 1'b0,  8'd26,  9'd279},{  1'b0, 1'b0,  8'd10,  9'd128},{  1'b0, 1'b0,   8'd4,  9'd154},{  1'b0, 1'b1,   8'd1,  9'd348},
{  1'b0, 1'b0, 8'd140,    9'd0},{  1'b0, 1'b0, 8'd139,    9'd0},{  1'b0, 1'b0,  8'd88,  9'd122},{  1'b0, 1'b0,  8'd68,    9'd0},{  1'b0, 1'b0,  8'd66,  9'd188},{  1'b0, 1'b0,  8'd32,  9'd223},{  1'b0, 1'b0,  8'd23,  9'd142},{  1'b0, 1'b0,  8'd22,  9'd135},{  1'b0, 1'b0,  8'd21,   9'd19},{  1'b0, 1'b0,   8'd7,  9'd197},{  1'b0, 1'b1,   8'd6,  9'd290},
{  1'b0, 1'b0, 8'd141,    9'd0},{  1'b0, 1'b0, 8'd140,    9'd0},{  1'b0, 1'b0,  8'd83,  9'd156},{  1'b0, 1'b0,  8'd69,    9'd0},{  1'b0, 1'b0,  8'd38,  9'd149},{  1'b0, 1'b0,  8'd30,  9'd335},{  1'b0, 1'b0,  8'd16,  9'd341},{  1'b0, 1'b0,  8'd14,  9'd333},{  1'b0, 1'b0,   8'd8,  9'd193},{  1'b0, 1'b0,   8'd3,  9'd327},{  1'b0, 1'b1,   8'd2,  9'd153},
{  1'b0, 1'b0, 8'd142,    9'd0},{  1'b0, 1'b0, 8'd141,    9'd0},{  1'b0, 1'b0, 8'd100,  9'd115},{  1'b0, 1'b0,  8'd70,    9'd0},{  1'b0, 1'b0,  8'd43,  9'd263},{  1'b0, 1'b0,  8'd23,  9'd238},{  1'b0, 1'b0,  8'd23,   9'd82},{  1'b0, 1'b0,  8'd19,  9'd184},{  1'b0, 1'b0,   8'd6,   9'd94},{  1'b0, 1'b0,   8'd3,   9'd72},{  1'b0, 1'b1,   8'd0,  9'd161},
{  1'b0, 1'b0, 8'd143,    9'd0},{  1'b0, 1'b0, 8'd142,    9'd0},{  1'b0, 1'b0,  8'd96,  9'd241},{  1'b0, 1'b0,  8'd71,    9'd0},{  1'b0, 1'b0,  8'd36,  9'd257},{  1'b0, 1'b0,  8'd27,  9'd324},{  1'b0, 1'b0,  8'd24,  9'd331},{  1'b0, 1'b0,  8'd13,  9'd164},{  1'b0, 1'b0,   8'd3,  9'd174},{  1'b0, 1'b0,   8'd3,  9'd160},{  1'b0, 1'b1,   8'd0,    9'd2},
{  1'b0, 1'b0, 8'd144,    9'd0},{  1'b0, 1'b0, 8'd143,    9'd0},{  1'b0, 1'b0, 8'd106,   9'd49},{  1'b0, 1'b0,  8'd72,    9'd0},{  1'b0, 1'b0,  8'd47,  9'd307},{  1'b0, 1'b0,  8'd26,  9'd293},{  1'b0, 1'b0,  8'd24,   9'd41},{  1'b0, 1'b0,  8'd13,   9'd10},{  1'b0, 1'b0,   8'd5,   9'd90},{  1'b0, 1'b0,   8'd4,   9'd15},{  1'b0, 1'b1,   8'd1,   9'd11},
{  1'b0, 1'b0, 8'd145,    9'd0},{  1'b0, 1'b0, 8'd144,    9'd0},{  1'b0, 1'b0, 8'd103,  9'd275},{  1'b0, 1'b0,  8'd73,    9'd0},{  1'b0, 1'b0,  8'd65,   9'd59},{  1'b0, 1'b0,  8'd24,  9'd101},{  1'b0, 1'b0,  8'd19,  9'd239},{  1'b0, 1'b0,  8'd17,  9'd335},{  1'b0, 1'b0,  8'd16,  9'd103},{  1'b0, 1'b0,   8'd5,  9'd208},{  1'b0, 1'b1,   8'd1,  9'd161},
{  1'b0, 1'b0, 8'd146,    9'd0},{  1'b0, 1'b0, 8'd145,    9'd0},{  1'b0, 1'b0,  8'd74,    9'd0},{  1'b0, 1'b0,  8'd74,   9'd68},{  1'b0, 1'b0,  8'd44,  9'd277},{  1'b0, 1'b0,  8'd35,  9'd192},{  1'b0, 1'b0,  8'd34,  9'd266},{  1'b0, 1'b0,  8'd25,  9'd324},{  1'b0, 1'b0,  8'd12,  9'd277},{  1'b0, 1'b0,  8'd11,  9'd253},{  1'b0, 1'b1,   8'd9,  9'd319},
{  1'b0, 1'b0, 8'd147,    9'd0},{  1'b0, 1'b0, 8'd146,    9'd0},{  1'b0, 1'b0,  8'd86,   9'd33},{  1'b0, 1'b0,  8'd75,    9'd0},{  1'b0, 1'b0,  8'd42,  9'd288},{  1'b0, 1'b0,  8'd30,   9'd55},{  1'b0, 1'b0,  8'd29,  9'd123},{  1'b0, 1'b0,  8'd22,  9'd119},{  1'b0, 1'b0,  8'd20,  9'd228},{  1'b0, 1'b0,  8'd20,  9'd303},{  1'b0, 1'b1,  8'd15,  9'd103},
{  1'b0, 1'b0, 8'd148,    9'd0},{  1'b0, 1'b0, 8'd147,    9'd0},{  1'b0, 1'b0, 8'd104,  9'd168},{  1'b0, 1'b0,  8'd76,    9'd0},{  1'b0, 1'b0,  8'd58,  9'd302},{  1'b0, 1'b0,  8'd26,   9'd98},{  1'b0, 1'b0,  8'd25,   9'd21},{  1'b0, 1'b0,  8'd20,  9'd213},{  1'b0, 1'b0,  8'd20,  9'd354},{  1'b0, 1'b0,  8'd15,   9'd15},{  1'b0, 1'b1,  8'd11,  9'd107},
{  1'b0, 1'b0, 8'd149,    9'd0},{  1'b0, 1'b0, 8'd148,    9'd0},{  1'b0, 1'b0,  8'd93,  9'd187},{  1'b0, 1'b0,  8'd77,    9'd0},{  1'b0, 1'b0,  8'd49,  9'd154},{  1'b0, 1'b0,  8'd34,  9'd346},{  1'b0, 1'b0,  8'd30,   9'd72},{  1'b0, 1'b0,  8'd25,  9'd267},{  1'b0, 1'b0,  8'd25,  9'd341},{  1'b0, 1'b0,   8'd9,   9'd40},{  1'b0, 1'b1,   8'd4,  9'd229},
{  1'b0, 1'b0, 8'd150,    9'd0},{  1'b0, 1'b0, 8'd149,    9'd0},{  1'b0, 1'b0,  8'd81,  9'd337},{  1'b0, 1'b0,  8'd78,    9'd0},{  1'b0, 1'b0,  8'd40,  9'd185},{  1'b0, 1'b0,  8'd31,  9'd288},{  1'b0, 1'b0,  8'd29,  9'd138},{  1'b0, 1'b0,  8'd22,  9'd327},{  1'b0, 1'b0,  8'd10,   9'd24},{  1'b0, 1'b0,   8'd2,  9'd157},{  1'b0, 1'b1,   8'd0,   9'd40},
{  1'b0, 1'b0, 8'd151,    9'd0},{  1'b0, 1'b0, 8'd150,    9'd0},{  1'b0, 1'b0,  8'd88,  9'd200},{  1'b0, 1'b0,  8'd79,    9'd0},{  1'b0, 1'b0,  8'd69,  9'd272},{  1'b0, 1'b0,  8'd34,  9'd156},{  1'b0, 1'b0,  8'd34,   9'd32},{  1'b0, 1'b0,  8'd24,  9'd181},{  1'b0, 1'b0,  8'd18,  9'd112},{  1'b0, 1'b0,  8'd12,   9'd16},{  1'b0, 1'b1,   8'd4,  9'd196},
{  1'b0, 1'b0, 8'd152,    9'd0},{  1'b0, 1'b0, 8'd151,    9'd0},{  1'b0, 1'b0,  8'd82,  9'd194},{  1'b0, 1'b0,  8'd80,    9'd0},{  1'b0, 1'b0,  8'd64,  9'd132},{  1'b0, 1'b0,  8'd26,  9'd273},{  1'b0, 1'b0,  8'd20,  9'd199},{  1'b0, 1'b0,  8'd15,  9'd350},{  1'b0, 1'b0,  8'd12,  9'd173},{  1'b0, 1'b0,   8'd8,  9'd298},{  1'b0, 1'b1,   8'd8,   9'd55},
{  1'b0, 1'b0, 8'd153,    9'd0},{  1'b0, 1'b0, 8'd152,    9'd0},{  1'b0, 1'b0, 8'd106,   9'd40},{  1'b0, 1'b0,  8'd81,    9'd0},{  1'b0, 1'b0,  8'd55,  9'd269},{  1'b0, 1'b0,  8'd33,  9'd118},{  1'b0, 1'b0,  8'd30,  9'd107},{  1'b0, 1'b0,  8'd30,  9'd311},{  1'b0, 1'b0,  8'd18,  9'd343},{  1'b0, 1'b0,   8'd9,   9'd78},{  1'b0, 1'b1,   8'd2,   9'd42},
{  1'b0, 1'b0, 8'd154,    9'd0},{  1'b0, 1'b0, 8'd153,    9'd0},{  1'b0, 1'b0,  8'd82,    9'd0},{  1'b0, 1'b0,  8'd77,  9'd104},{  1'b0, 1'b0,  8'd65,  9'd243},{  1'b0, 1'b0,  8'd34,   9'd99},{  1'b0, 1'b0,  8'd33,   9'd89},{  1'b0, 1'b0,  8'd24,  9'd182},{  1'b0, 1'b0,  8'd24,  9'd332},{  1'b0, 1'b0,   8'd8,  9'd344},{  1'b0, 1'b1,   8'd8,   9'd30},
{  1'b0, 1'b0, 8'd155,    9'd0},{  1'b0, 1'b0, 8'd154,    9'd0},{  1'b0, 1'b0,  8'd91,   9'd56},{  1'b0, 1'b0,  8'd83,    9'd0},{  1'b0, 1'b0,  8'd54,  9'd274},{  1'b0, 1'b0,  8'd35,   9'd39},{  1'b0, 1'b0,  8'd26,  9'd261},{  1'b0, 1'b0,  8'd26,   9'd78},{  1'b0, 1'b0,  8'd21,  9'd324},{  1'b0, 1'b0,  8'd13,   9'd50},{  1'b0, 1'b1,   8'd7,  9'd125},
{  1'b0, 1'b0, 8'd156,    9'd0},{  1'b0, 1'b0, 8'd155,    9'd0},{  1'b0, 1'b0,  8'd84,    9'd0},{  1'b0, 1'b0,  8'd72,  9'd193},{  1'b0, 1'b0,  8'd71,  9'd240},{  1'b0, 1'b0,  8'd27,  9'd310},{  1'b0, 1'b0,  8'd21,  9'd179},{  1'b0, 1'b0,  8'd21,  9'd354},{  1'b0, 1'b0,  8'd13,  9'd318},{  1'b0, 1'b0,  8'd12,  9'd262},{  1'b0, 1'b1,   8'd4,  9'd291},
{  1'b0, 1'b0, 8'd157,    9'd0},{  1'b0, 1'b0, 8'd156,    9'd0},{  1'b0, 1'b0,  8'd85,    9'd0},{  1'b0, 1'b0,  8'd73,  9'd312},{  1'b0, 1'b0,  8'd56,   9'd50},{  1'b0, 1'b0,  8'd28,   9'd56},{  1'b0, 1'b0,  8'd23,  9'd247},{  1'b0, 1'b0,  8'd20,   9'd24},{  1'b0, 1'b0,  8'd13,  9'd179},{  1'b0, 1'b0,   8'd9,  9'd274},{  1'b0, 1'b1,   8'd3,  9'd308},
{  1'b0, 1'b0, 8'd158,    9'd0},{  1'b0, 1'b0, 8'd157,    9'd0},{  1'b0, 1'b0, 8'd107,   9'd47},{  1'b0, 1'b0,  8'd86,    9'd0},{  1'b0, 1'b0,  8'd37,   9'd41},{  1'b0, 1'b0,  8'd32,  9'd137},{  1'b0, 1'b0,  8'd29,  9'd327},{  1'b0, 1'b0,  8'd20,  9'd252},{  1'b0, 1'b0,  8'd14,   9'd11},{  1'b0, 1'b0,   8'd7,  9'd233},{  1'b0, 1'b1,   8'd5,  9'd131},
{  1'b0, 1'b0, 8'd159,    9'd0},{  1'b0, 1'b0, 8'd158,    9'd0},{  1'b0, 1'b0,  8'd87,    9'd0},{  1'b0, 1'b0,  8'd84,  9'd215},{  1'b0, 1'b0,  8'd57,  9'd185},{  1'b0, 1'b0,  8'd34,  9'd344},{  1'b0, 1'b0,  8'd33,  9'd264},{  1'b0, 1'b0,  8'd23,   9'd75},{  1'b0, 1'b0,  8'd14,   9'd69},{  1'b0, 1'b0,  8'd12,  9'd278},{  1'b0, 1'b1,   8'd1,  9'd312},
{  1'b0, 1'b0, 8'd160,    9'd0},{  1'b0, 1'b0, 8'd159,    9'd0},{  1'b0, 1'b0,  8'd88,    9'd0},{  1'b0, 1'b0,  8'd87,  9'd346},{  1'b0, 1'b0,  8'd39,  9'd108},{  1'b0, 1'b0,  8'd33,  9'd145},{  1'b0, 1'b0,  8'd23,  9'd223},{  1'b0, 1'b0,  8'd21,  9'd117},{  1'b0, 1'b0,  8'd21,   9'd56},{  1'b0, 1'b0,  8'd14,  9'd122},{  1'b0, 1'b1,   8'd7,   9'd76},
{  1'b0, 1'b0, 8'd161,    9'd0},{  1'b0, 1'b0, 8'd160,    9'd0},{  1'b0, 1'b0,  8'd89,    9'd0},{  1'b0, 1'b0,  8'd78,  9'd177},{  1'b0, 1'b0,  8'd61,   9'd51},{  1'b0, 1'b0,  8'd28,   9'd68},{  1'b0, 1'b0,  8'd13,  9'd114},{  1'b0, 1'b0,   8'd9,  9'd312},{  1'b0, 1'b0,   8'd9,   9'd33},{  1'b0, 1'b0,   8'd7,  9'd330},{  1'b0, 1'b1,   8'd0,  9'd277},
{  1'b0, 1'b0, 8'd162,    9'd0},{  1'b0, 1'b0, 8'd161,    9'd0},{  1'b0, 1'b0, 8'd105,  9'd107},{  1'b0, 1'b0,  8'd90,    9'd0},{  1'b0, 1'b0,  8'd68,  9'd322},{  1'b0, 1'b0,  8'd32,   9'd35},{  1'b0, 1'b0,  8'd19,  9'd351},{  1'b0, 1'b0,  8'd17,   9'd51},{  1'b0, 1'b0,  8'd16,  9'd128},{  1'b0, 1'b0,  8'd16,  9'd229},{  1'b0, 1'b1,  8'd16,  9'd203},
{  1'b0, 1'b0, 8'd163,    9'd0},{  1'b0, 1'b0, 8'd162,    9'd0},{  1'b0, 1'b0, 8'd101,  9'd278},{  1'b0, 1'b0,  8'd91,    9'd0},{  1'b0, 1'b0,  8'd63,   9'd79},{  1'b0, 1'b0,  8'd31,  9'd164},{  1'b0, 1'b0,  8'd29,  9'd183},{  1'b0, 1'b0,  8'd27,  9'd111},{  1'b0, 1'b0,  8'd18,  9'd230},{  1'b0, 1'b0,  8'd12,  9'd291},{  1'b0, 1'b1,   8'd1,   9'd89},
{  1'b0, 1'b0, 8'd164,    9'd0},{  1'b0, 1'b0, 8'd163,    9'd0},{  1'b0, 1'b0, 8'd105,  9'd316},{  1'b0, 1'b0,  8'd92,    9'd0},{  1'b0, 1'b0,  8'd68,  9'd161},{  1'b0, 1'b0,  8'd22,    9'd1},{  1'b0, 1'b0,  8'd22,   9'd25},{  1'b0, 1'b0,  8'd18,  9'd345},{  1'b0, 1'b0,  8'd18,  9'd359},{  1'b0, 1'b0,  8'd16,   9'd50},{  1'b0, 1'b1,  8'd15,   9'd65},
{  1'b0, 1'b0, 8'd165,    9'd0},{  1'b0, 1'b0, 8'd164,    9'd0},{  1'b0, 1'b0,  8'd93,    9'd0},{  1'b0, 1'b0,  8'd85,  9'd130},{  1'b0, 1'b0,  8'd61,   9'd88},{  1'b0, 1'b0,  8'd34,  9'd100},{  1'b0, 1'b0,  8'd19,   9'd51},{  1'b0, 1'b0,  8'd16,  9'd219},{  1'b0, 1'b0,  8'd12,   9'd85},{  1'b0, 1'b0,   8'd9,  9'd264},{  1'b0, 1'b1,   8'd2,  9'd239},
{  1'b0, 1'b0, 8'd166,    9'd0},{  1'b0, 1'b0, 8'd165,    9'd0},{  1'b0, 1'b0,  8'd95,   9'd21},{  1'b0, 1'b0,  8'd94,    9'd0},{  1'b0, 1'b0,  8'd67,   9'd24},{  1'b0, 1'b0,  8'd34,   9'd40},{  1'b0, 1'b0,  8'd31,  9'd110},{  1'b0, 1'b0,  8'd28,  9'd100},{  1'b0, 1'b0,  8'd25,  9'd244},{  1'b0, 1'b0,   8'd5,   9'd14},{  1'b0, 1'b1,   8'd0,  9'd142},
{  1'b0, 1'b0, 8'd167,    9'd0},{  1'b0, 1'b0, 8'd166,    9'd0},{  1'b0, 1'b0,  8'd95,    9'd0},{  1'b0, 1'b0,  8'd74,  9'd174},{  1'b0, 1'b0,  8'd39,  9'd170},{  1'b0, 1'b0,  8'd19,   9'd70},{  1'b0, 1'b0,  8'd16,  9'd329},{  1'b0, 1'b0,  8'd12,  9'd332},{  1'b0, 1'b0,   8'd5,  9'd197},{  1'b0, 1'b0,   8'd4,  9'd148},{  1'b0, 1'b1,   8'd3,  9'd352},
{  1'b0, 1'b0, 8'd168,    9'd0},{  1'b0, 1'b0, 8'd167,    9'd0},{  1'b0, 1'b0,  8'd96,    9'd0},{  1'b0, 1'b0,  8'd80,   9'd15},{  1'b0, 1'b0,  8'd71,  9'd190},{  1'b0, 1'b0,  8'd35,  9'd208},{  1'b0, 1'b0,  8'd33,  9'd158},{  1'b0, 1'b0,  8'd28,   9'd97},{  1'b0, 1'b0,  8'd25,  9'd250},{  1'b0, 1'b0,   8'd6,  9'd308},{  1'b0, 1'b1,   8'd2,  9'd199},
{  1'b0, 1'b0, 8'd169,    9'd0},{  1'b0, 1'b0, 8'd168,    9'd0},{  1'b0, 1'b0, 8'd100,   9'd18},{  1'b0, 1'b0,  8'd97,    9'd0},{  1'b0, 1'b0,  8'd50,  9'd191},{  1'b0, 1'b0,  8'd21,  9'd309},{  1'b0, 1'b0,  8'd20,  9'd173},{  1'b0, 1'b0,  8'd18,  9'd282},{  1'b0, 1'b0,  8'd14,  9'd337},{  1'b0, 1'b0,   8'd5,  9'd231},{  1'b0, 1'b1,   8'd3,  9'd273},
{  1'b0, 1'b0, 8'd170,    9'd0},{  1'b0, 1'b0, 8'd169,    9'd0},{  1'b0, 1'b0,  8'd98,    9'd0},{  1'b0, 1'b0,  8'd84,   9'd64},{  1'b0, 1'b0,  8'd37,  9'd145},{  1'b0, 1'b0,  8'd33,  9'd227},{  1'b0, 1'b0,  8'd32,  9'd156},{  1'b0, 1'b0,  8'd30,  9'd184},{  1'b0, 1'b0,  8'd29,  9'd296},{  1'b0, 1'b0,  8'd12,   9'd60},{  1'b0, 1'b1,   8'd0,  9'd114},
{  1'b0, 1'b0, 8'd171,    9'd0},{  1'b0, 1'b0, 8'd170,    9'd0},{  1'b0, 1'b0,  8'd99,    9'd0},{  1'b0, 1'b0,  8'd73,   9'd92},{  1'b0, 1'b0,  8'd66,  9'd313},{  1'b0, 1'b0,  8'd32,  9'd316},{  1'b0, 1'b0,  8'd31,  9'd357},{  1'b0, 1'b0,  8'd28,  9'd339},{  1'b0, 1'b0,  8'd22,  9'd348},{  1'b0, 1'b0,   8'd4,   9'd78},{  1'b0, 1'b1,   8'd1,  9'd313},
{  1'b0, 1'b0, 8'd172,    9'd0},{  1'b0, 1'b0, 8'd171,    9'd0},{  1'b0, 1'b0, 8'd100,    9'd0},{  1'b0, 1'b0,  8'd78,  9'd338},{  1'b0, 1'b0,  8'd45,  9'd156},{  1'b0, 1'b0,  8'd35,  9'd321},{  1'b0, 1'b0,  8'd34,  9'd225},{  1'b0, 1'b0,  8'd23,  9'd293},{  1'b0, 1'b0,  8'd10,  9'd152},{  1'b0, 1'b0,   8'd8,  9'd229},{  1'b0, 1'b1,   8'd6,   9'd95},
{  1'b0, 1'b0, 8'd173,    9'd0},{  1'b0, 1'b0, 8'd172,    9'd0},{  1'b0, 1'b0, 8'd107,  9'd107},{  1'b0, 1'b0, 8'd101,    9'd0},{  1'b0, 1'b0,  8'd70,  9'd188},{  1'b0, 1'b0,  8'd35,   9'd82},{  1'b0, 1'b0,  8'd31,  9'd236},{  1'b0, 1'b0,  8'd26,  9'd194},{  1'b0, 1'b0,  8'd17,  9'd235},{  1'b0, 1'b0,  8'd14,  9'd153},{  1'b0, 1'b1,   8'd7,  9'd273},
{  1'b0, 1'b0, 8'd174,    9'd0},{  1'b0, 1'b0, 8'd173,    9'd0},{  1'b0, 1'b0, 8'd102,    9'd0},{  1'b0, 1'b0,  8'd87,  9'd342},{  1'b0, 1'b0,  8'd70,  9'd186},{  1'b0, 1'b0,  8'd29,  9'd196},{  1'b0, 1'b0,  8'd24,  9'd340},{  1'b0, 1'b0,  8'd21,   9'd88},{  1'b0, 1'b0,  8'd20,  9'd242},{  1'b0, 1'b0,  8'd19,  9'd341},{  1'b0, 1'b1,   8'd5,   9'd19},
{  1'b0, 1'b0, 8'd175,    9'd0},{  1'b0, 1'b0, 8'd174,    9'd0},{  1'b0, 1'b0, 8'd103,    9'd0},{  1'b0, 1'b0,  8'd89,   9'd17},{  1'b0, 1'b0,  8'd46,  9'd286},{  1'b0, 1'b0,  8'd34,  9'd175},{  1'b0, 1'b0,  8'd33,   9'd79},{  1'b0, 1'b0,  8'd28,  9'd147},{  1'b0, 1'b0,  8'd10,   9'd37},{  1'b0, 1'b0,   8'd6,  9'd217},{  1'b0, 1'b1,   8'd6,  9'd299},
{  1'b0, 1'b0, 8'd176,    9'd0},{  1'b0, 1'b0, 8'd175,    9'd0},{  1'b0, 1'b0, 8'd104,    9'd0},{  1'b0, 1'b0,  8'd95,   9'd83},{  1'b0, 1'b0,  8'd53,   9'd80},{  1'b0, 1'b0,  8'd26,  9'd173},{  1'b0, 1'b0,  8'd17,  9'd315},{  1'b0, 1'b0,  8'd14,  9'd111},{  1'b0, 1'b0,   8'd6,    9'd6},{  1'b0, 1'b0,   8'd5,  9'd119},{  1'b0, 1'b1,   8'd4,  9'd216},
{  1'b0, 1'b0, 8'd177,    9'd0},{  1'b0, 1'b0, 8'd176,    9'd0},{  1'b0, 1'b0, 8'd105,    9'd0},{  1'b0, 1'b0,  8'd93,   9'd84},{  1'b0, 1'b0,  8'd48,  9'd305},{  1'b0, 1'b0,  8'd35,    9'd7},{  1'b0, 1'b0,  8'd28,  9'd198},{  1'b0, 1'b0,  8'd19,  9'd284},{  1'b0, 1'b0,  8'd18,  9'd186},{  1'b0, 1'b0,  8'd12,  9'd344},{  1'b0, 1'b1,  8'd11,  9'd353},
{  1'b0, 1'b0, 8'd178,    9'd0},{  1'b0, 1'b0, 8'd177,    9'd0},{  1'b0, 1'b0, 8'd106,    9'd0},{  1'b0, 1'b0,  8'd90,  9'd288},{  1'b0, 1'b0,  8'd46,  9'd208},{  1'b0, 1'b0,  8'd28,   9'd14},{  1'b0, 1'b0,  8'd28,   9'd59},{  1'b0, 1'b0,  8'd24,  9'd274},{  1'b0, 1'b0,  8'd19,  9'd136},{  1'b0, 1'b0,  8'd16,  9'd311},{  1'b0, 1'b1,  8'd13,  9'd154},
{  1'b0, 1'b0, 8'd179,    9'd0},{  1'b0, 1'b0, 8'd178,    9'd0},{  1'b0, 1'b0, 8'd107,    9'd0},{  1'b0, 1'b0,  8'd98,  9'd285},{  1'b0, 1'b0,  8'd54,   9'd58},{  1'b0, 1'b0,  8'd31,  9'd341},{  1'b0, 1'b0,  8'd21,  9'd112},{  1'b0, 1'b0,  8'd21,  9'd289},{  1'b0, 1'b0,  8'd19,  9'd196},{  1'b0, 1'b0,  8'd15,   9'd76},{  1'b0, 1'b1,  8'd10,   9'd10}
};
localparam bit [18 : 0] cLARGE_HS_V_TAB_3BY5_PACKED[cLARGE_HS_TAB_3BY5_PACKED_SIZE] = '{
{8'd179, 1'b0,   10'd0},{8'd179, 1'b1, 10'd781},
{8'd178, 1'b0, 10'd770},{8'd178, 1'b1, 10'd782},
{8'd177, 1'b0, 10'd759},{8'd177, 1'b1, 10'd771},
{8'd176, 1'b0, 10'd748},{8'd176, 1'b1, 10'd760},
{8'd175, 1'b0, 10'd737},{8'd175, 1'b1, 10'd749},
{8'd174, 1'b0, 10'd726},{8'd174, 1'b1, 10'd738},
{8'd173, 1'b0, 10'd715},{8'd173, 1'b1, 10'd727},
{8'd172, 1'b0, 10'd704},{8'd172, 1'b1, 10'd716},
{8'd171, 1'b0, 10'd693},{8'd171, 1'b1, 10'd705},
{8'd170, 1'b0, 10'd682},{8'd170, 1'b1, 10'd694},
{8'd169, 1'b0, 10'd671},{8'd169, 1'b1, 10'd683},
{8'd168, 1'b0, 10'd660},{8'd168, 1'b1, 10'd672},
{8'd167, 1'b0, 10'd649},{8'd167, 1'b1, 10'd661},
{8'd166, 1'b0, 10'd638},{8'd166, 1'b1, 10'd650},
{8'd165, 1'b0, 10'd627},{8'd165, 1'b1, 10'd639},
{8'd164, 1'b0, 10'd616},{8'd164, 1'b1, 10'd628},
{8'd163, 1'b0, 10'd605},{8'd163, 1'b1, 10'd617},
{8'd162, 1'b0, 10'd594},{8'd162, 1'b1, 10'd606},
{8'd161, 1'b0, 10'd583},{8'd161, 1'b1, 10'd595},
{8'd160, 1'b0, 10'd572},{8'd160, 1'b1, 10'd584},
{8'd159, 1'b0, 10'd561},{8'd159, 1'b1, 10'd573},
{8'd158, 1'b0, 10'd550},{8'd158, 1'b1, 10'd562},
{8'd157, 1'b0, 10'd539},{8'd157, 1'b1, 10'd551},
{8'd156, 1'b0, 10'd528},{8'd156, 1'b1, 10'd540},
{8'd155, 1'b0, 10'd517},{8'd155, 1'b1, 10'd529},
{8'd154, 1'b0, 10'd506},{8'd154, 1'b1, 10'd518},
{8'd153, 1'b0, 10'd495},{8'd153, 1'b1, 10'd507},
{8'd152, 1'b0, 10'd484},{8'd152, 1'b1, 10'd496},
{8'd151, 1'b0, 10'd473},{8'd151, 1'b1, 10'd485},
{8'd150, 1'b0, 10'd462},{8'd150, 1'b1, 10'd474},
{8'd149, 1'b0, 10'd451},{8'd149, 1'b1, 10'd463},
{8'd148, 1'b0, 10'd440},{8'd148, 1'b1, 10'd452},
{8'd147, 1'b0, 10'd429},{8'd147, 1'b1, 10'd441},
{8'd146, 1'b0, 10'd418},{8'd146, 1'b1, 10'd430},
{8'd145, 1'b0, 10'd407},{8'd145, 1'b1, 10'd419},
{8'd144, 1'b0, 10'd396},{8'd144, 1'b1, 10'd408},
{8'd143, 1'b0, 10'd385},{8'd143, 1'b1, 10'd397},
{8'd142, 1'b0, 10'd374},{8'd142, 1'b1, 10'd386},
{8'd141, 1'b0, 10'd363},{8'd141, 1'b1, 10'd375},
{8'd140, 1'b0, 10'd352},{8'd140, 1'b1, 10'd364},
{8'd139, 1'b0, 10'd341},{8'd139, 1'b1, 10'd353},
{8'd138, 1'b0, 10'd330},{8'd138, 1'b1, 10'd342},
{8'd137, 1'b0, 10'd319},{8'd137, 1'b1, 10'd331},
{8'd136, 1'b0, 10'd308},{8'd136, 1'b1, 10'd320},
{8'd135, 1'b0, 10'd297},{8'd135, 1'b1, 10'd309},
{8'd134, 1'b0, 10'd286},{8'd134, 1'b1, 10'd298},
{8'd133, 1'b0, 10'd275},{8'd133, 1'b1, 10'd287},
{8'd132, 1'b0, 10'd264},{8'd132, 1'b1, 10'd276},
{8'd131, 1'b0, 10'd253},{8'd131, 1'b1, 10'd265},
{8'd130, 1'b0, 10'd242},{8'd130, 1'b1, 10'd254},
{8'd129, 1'b0, 10'd231},{8'd129, 1'b1, 10'd243},
{8'd128, 1'b0, 10'd220},{8'd128, 1'b1, 10'd232},
{8'd127, 1'b0, 10'd209},{8'd127, 1'b1, 10'd221},
{8'd126, 1'b0, 10'd198},{8'd126, 1'b1, 10'd210},
{8'd125, 1'b0, 10'd187},{8'd125, 1'b1, 10'd199},
{8'd124, 1'b0, 10'd176},{8'd124, 1'b1, 10'd188},
{8'd123, 1'b0, 10'd165},{8'd123, 1'b1, 10'd177},
{8'd122, 1'b0, 10'd154},{8'd122, 1'b1, 10'd166},
{8'd121, 1'b0, 10'd143},{8'd121, 1'b1, 10'd155},
{8'd120, 1'b0, 10'd132},{8'd120, 1'b1, 10'd144},
{8'd119, 1'b0, 10'd121},{8'd119, 1'b1, 10'd133},
{8'd118, 1'b0, 10'd110},{8'd118, 1'b1, 10'd122},
{8'd117, 1'b0,  10'd99},{8'd117, 1'b1, 10'd111},
{8'd116, 1'b0,  10'd88},{8'd116, 1'b1, 10'd100},
{8'd115, 1'b0,  10'd77},{8'd115, 1'b1,  10'd89},
{8'd114, 1'b0,  10'd66},{8'd114, 1'b1,  10'd78},
{8'd113, 1'b0,  10'd55},{8'd113, 1'b1,  10'd67},
{8'd112, 1'b0,  10'd44},{8'd112, 1'b1,  10'd56},
{8'd111, 1'b0,  10'd33},{8'd111, 1'b1,  10'd45},
{8'd110, 1'b0,  10'd22},{8'd110, 1'b1,  10'd34},
{8'd109, 1'b0,  10'd11},{8'd109, 1'b1,  10'd23},
{8'd108, 1'b0,   10'd1},{8'd108, 1'b1,  10'd12},
{8'd107, 1'b0, 10'd552},{8'd107, 1'b0, 10'd717},{8'd107, 1'b1, 10'd783},
{8'd106, 1'b0, 10'd398},{8'd106, 1'b0, 10'd497},{8'd106, 1'b1, 10'd772},
{8'd105, 1'b0, 10'd596},{8'd105, 1'b0, 10'd618},{8'd105, 1'b1, 10'd761},
{8'd104, 1'b0,  10'd35},{8'd104, 1'b0, 10'd442},{8'd104, 1'b1, 10'd750},
{8'd103, 1'b0, 10'd112},{8'd103, 1'b0, 10'd409},{8'd103, 1'b1, 10'd739},
{8'd102, 1'b0, 10'd178},{8'd102, 1'b0, 10'd244},{8'd102, 1'b1, 10'd728},
{8'd101, 1'b0,   10'd2},{8'd101, 1'b0, 10'd607},{8'd101, 1'b1, 10'd718},
{8'd100, 1'b0, 10'd376},{8'd100, 1'b0, 10'd673},{8'd100, 1'b1, 10'd706},
{ 8'd99, 1'b0, 10'd200},{ 8'd99, 1'b0, 10'd332},{ 8'd99, 1'b1, 10'd695},
{ 8'd98, 1'b0,  10'd68},{ 8'd98, 1'b0, 10'd684},{ 8'd98, 1'b1, 10'd784},
{ 8'd97, 1'b0,  10'd13},{ 8'd97, 1'b0,  10'd79},{ 8'd97, 1'b1, 10'd674},
{ 8'd96, 1'b0,  10'd46},{ 8'd96, 1'b0, 10'd387},{ 8'd96, 1'b1, 10'd662},
{ 8'd95, 1'b0, 10'd640},{ 8'd95, 1'b0, 10'd651},{ 8'd95, 1'b1, 10'd751},
{ 8'd94, 1'b0,  10'd57},{ 8'd94, 1'b0, 10'd134},{ 8'd94, 1'b1, 10'd641},
{ 8'd93, 1'b0, 10'd453},{ 8'd93, 1'b0, 10'd629},{ 8'd93, 1'b1, 10'd762},
{ 8'd92, 1'b0,  10'd24},{ 8'd92, 1'b0, 10'd222},{ 8'd92, 1'b1, 10'd619},
{ 8'd91, 1'b0, 10'd211},{ 8'd91, 1'b0, 10'd519},{ 8'd91, 1'b1, 10'd608},
{ 8'd90, 1'b0, 10'd189},{ 8'd90, 1'b0, 10'd597},{ 8'd90, 1'b1, 10'd773},
{ 8'd89, 1'b0, 10'd156},{ 8'd89, 1'b0, 10'd585},{ 8'd89, 1'b1, 10'd740},
{ 8'd88, 1'b0, 10'd354},{ 8'd88, 1'b0, 10'd475},{ 8'd88, 1'b1, 10'd574},
{ 8'd87, 1'b0, 10'd563},{ 8'd87, 1'b0, 10'd575},{ 8'd87, 1'b1, 10'd729},
{ 8'd86, 1'b0, 10'd266},{ 8'd86, 1'b0, 10'd431},{ 8'd86, 1'b1, 10'd553},
{ 8'd85, 1'b0, 10'd343},{ 8'd85, 1'b0, 10'd541},{ 8'd85, 1'b1, 10'd630},
{ 8'd84, 1'b0, 10'd530},{ 8'd84, 1'b0, 10'd564},{ 8'd84, 1'b1, 10'd685},
{ 8'd83, 1'b0, 10'd299},{ 8'd83, 1'b0, 10'd365},{ 8'd83, 1'b1, 10'd520},
{ 8'd82, 1'b0, 10'd123},{ 8'd82, 1'b0, 10'd486},{ 8'd82, 1'b1, 10'd508},
{ 8'd81, 1'b0, 10'd145},{ 8'd81, 1'b0, 10'd464},{ 8'd81, 1'b1, 10'd498},
{ 8'd80, 1'b0, 10'd167},{ 8'd80, 1'b0, 10'd487},{ 8'd80, 1'b1, 10'd663},
{ 8'd79, 1'b0,  10'd90},{ 8'd79, 1'b0, 10'd255},{ 8'd79, 1'b1, 10'd476},
{ 8'd78, 1'b0, 10'd465},{ 8'd78, 1'b0, 10'd586},{ 8'd78, 1'b1, 10'd707},
{ 8'd77, 1'b0, 10'd101},{ 8'd77, 1'b0, 10'd454},{ 8'd77, 1'b1, 10'd509},
{ 8'd76, 1'b0, 10'd277},{ 8'd76, 1'b0, 10'd288},{ 8'd76, 1'b1, 10'd443},
{ 8'd75, 1'b0, 10'd233},{ 8'd75, 1'b0, 10'd321},{ 8'd75, 1'b1, 10'd432},
{ 8'd74, 1'b0, 10'd420},{ 8'd74, 1'b0, 10'd421},{ 8'd74, 1'b1, 10'd652},
{ 8'd73, 1'b0, 10'd410},{ 8'd73, 1'b0, 10'd542},{ 8'd73, 1'b1, 10'd696},
{ 8'd72, 1'b0, 10'd310},{ 8'd72, 1'b0, 10'd399},{ 8'd72, 1'b1, 10'd531},
{ 8'd71, 1'b0, 10'd388},{ 8'd71, 1'b0, 10'd532},{ 8'd71, 1'b1, 10'd664},
{ 8'd70, 1'b0, 10'd377},{ 8'd70, 1'b0, 10'd719},{ 8'd70, 1'b1, 10'd730},
{ 8'd69, 1'b0, 10'd157},{ 8'd69, 1'b0, 10'd366},{ 8'd69, 1'b1, 10'd477},
{ 8'd68, 1'b0, 10'd355},{ 8'd68, 1'b0, 10'd598},{ 8'd68, 1'b1, 10'd620},
{ 8'd67, 1'b0, 10'd102},{ 8'd67, 1'b0, 10'd344},{ 8'd67, 1'b1, 10'd642},
{ 8'd66, 1'b0, 10'd333},{ 8'd66, 1'b0, 10'd356},{ 8'd66, 1'b1, 10'd697},
{ 8'd65, 1'b0, 10'd322},{ 8'd65, 1'b0, 10'd411},{ 8'd65, 1'b1, 10'd510},
{ 8'd64, 1'b0,  10'd25},{ 8'd64, 1'b0, 10'd311},{ 8'd64, 1'b1, 10'd488},
{ 8'd63, 1'b0, 10'd223},{ 8'd63, 1'b0, 10'd300},{ 8'd63, 1'b1, 10'd609},
{ 8'd62, 1'b0, 10'd234},{ 8'd62, 1'b0, 10'd267},{ 8'd62, 1'b1, 10'd289},
{ 8'd61, 1'b0, 10'd278},{ 8'd61, 1'b0, 10'd587},{ 8'd61, 1'b1, 10'd631},
{ 8'd60, 1'b0, 10'd168},{ 8'd60, 1'b0, 10'd190},{ 8'd60, 1'b1, 10'd268},
{ 8'd59, 1'b0, 10'd212},{ 8'd59, 1'b0, 10'd256},{ 8'd59, 1'b1, 10'd323},
{ 8'd58, 1'b0, 10'd201},{ 8'd58, 1'b0, 10'd245},{ 8'd58, 1'b1, 10'd444},
{ 8'd57, 1'b0,  10'd36},{ 8'd57, 1'b0, 10'd235},{ 8'd57, 1'b1, 10'd565},
{ 8'd56, 1'b0, 10'd124},{ 8'd56, 1'b0, 10'd224},{ 8'd56, 1'b1, 10'd543},
{ 8'd55, 1'b0,  10'd47},{ 8'd55, 1'b0, 10'd213},{ 8'd55, 1'b1, 10'd499},
{ 8'd54, 1'b0, 10'd202},{ 8'd54, 1'b0, 10'd521},{ 8'd54, 1'b1, 10'd785},
{ 8'd53, 1'b0, 10'd191},{ 8'd53, 1'b0, 10'd334},{ 8'd53, 1'b1, 10'd752},
{ 8'd52, 1'b0, 10'd179},{ 8'd52, 1'b0, 10'd290},{ 8'd52, 1'b1, 10'd345},
{ 8'd51, 1'b0, 10'd113},{ 8'd51, 1'b0, 10'd169},{ 8'd51, 1'b1, 10'd279},
{ 8'd50, 1'b0,  10'd69},{ 8'd50, 1'b0, 10'd158},{ 8'd50, 1'b1, 10'd675},
{ 8'd49, 1'b0, 10'd146},{ 8'd49, 1'b0, 10'd246},{ 8'd49, 1'b1, 10'd455},
{ 8'd48, 1'b0,  10'd58},{ 8'd48, 1'b0, 10'd135},{ 8'd48, 1'b1, 10'd763},
{ 8'd47, 1'b0, 10'd125},{ 8'd47, 1'b0, 10'd312},{ 8'd47, 1'b1, 10'd400},
{ 8'd46, 1'b0, 10'd114},{ 8'd46, 1'b0, 10'd741},{ 8'd46, 1'b1, 10'd774},
{ 8'd45, 1'b0,  10'd80},{ 8'd45, 1'b0, 10'd103},{ 8'd45, 1'b1, 10'd708},
{ 8'd44, 1'b0,  10'd14},{ 8'd44, 1'b0,  10'd91},{ 8'd44, 1'b1, 10'd422},
{ 8'd43, 1'b0,  10'd81},{ 8'd43, 1'b0, 10'd301},{ 8'd43, 1'b1, 10'd378},
{ 8'd42, 1'b0,  10'd70},{ 8'd42, 1'b0, 10'd257},{ 8'd42, 1'b1, 10'd433},
{ 8'd41, 1'b0,  10'd59},{ 8'd41, 1'b0, 10'd136},{ 8'd41, 1'b1, 10'd180},
{ 8'd40, 1'b0,   10'd3},{ 8'd40, 1'b0,  10'd48},{ 8'd40, 1'b1, 10'd466},
{ 8'd39, 1'b0,  10'd37},{ 8'd39, 1'b0, 10'd576},{ 8'd39, 1'b1, 10'd653},
{ 8'd38, 1'b0,  10'd26},{ 8'd38, 1'b0,  10'd92},{ 8'd38, 1'b1, 10'd367},
{ 8'd37, 1'b0,  10'd15},{ 8'd37, 1'b0, 10'd554},{ 8'd37, 1'b1, 10'd686},
{ 8'd36, 1'b0,   10'd4},{ 8'd36, 1'b0, 10'd147},{ 8'd36, 1'b1, 10'd389},
{ 8'd35, 1'b0,  10'd93},{ 8'd35, 1'b0, 10'd137},{ 8'd35, 1'b0, 10'd192},{ 8'd35, 1'b0, 10'd269},{ 8'd35, 1'b0, 10'd291},{ 8'd35, 1'b0, 10'd302},{ 8'd35, 1'b0, 10'd423},{ 8'd35, 1'b0, 10'd522},{ 8'd35, 1'b0, 10'd665},{ 8'd35, 1'b0, 10'd709},{ 8'd35, 1'b0, 10'd720},{ 8'd35, 1'b1, 10'd764},
{ 8'd34, 1'b0,  10'd27},{ 8'd34, 1'b0, 10'd148},{ 8'd34, 1'b0, 10'd424},{ 8'd34, 1'b0, 10'd456},{ 8'd34, 1'b0, 10'd478},{ 8'd34, 1'b0, 10'd479},{ 8'd34, 1'b0, 10'd511},{ 8'd34, 1'b0, 10'd566},{ 8'd34, 1'b0, 10'd632},{ 8'd34, 1'b0, 10'd643},{ 8'd34, 1'b0, 10'd710},{ 8'd34, 1'b1, 10'd742},
{ 8'd33, 1'b0,   10'd5},{ 8'd33, 1'b0,  10'd16},{ 8'd33, 1'b0,  10'd28},{ 8'd33, 1'b0, 10'd138},{ 8'd33, 1'b0, 10'd346},{ 8'd33, 1'b0, 10'd500},{ 8'd33, 1'b0, 10'd512},{ 8'd33, 1'b0, 10'd567},{ 8'd33, 1'b0, 10'd577},{ 8'd33, 1'b0, 10'd666},{ 8'd33, 1'b0, 10'd687},{ 8'd33, 1'b1, 10'd743},
{ 8'd32, 1'b0,   10'd6},{ 8'd32, 1'b0, 10'd170},{ 8'd32, 1'b0, 10'd225},{ 8'd32, 1'b0, 10'd280},{ 8'd32, 1'b0, 10'd303},{ 8'd32, 1'b0, 10'd313},{ 8'd32, 1'b0, 10'd347},{ 8'd32, 1'b0, 10'd357},{ 8'd32, 1'b0, 10'd555},{ 8'd32, 1'b0, 10'd599},{ 8'd32, 1'b0, 10'd688},{ 8'd32, 1'b1, 10'd698},
{ 8'd31, 1'b0,  10'd60},{ 8'd31, 1'b0,  10'd82},{ 8'd31, 1'b0, 10'd104},{ 8'd31, 1'b0, 10'd149},{ 8'd31, 1'b0, 10'd171},{ 8'd31, 1'b0, 10'd214},{ 8'd31, 1'b0, 10'd467},{ 8'd31, 1'b0, 10'd610},{ 8'd31, 1'b0, 10'd644},{ 8'd31, 1'b0, 10'd699},{ 8'd31, 1'b0, 10'd721},{ 8'd31, 1'b1, 10'd786},
{ 8'd30, 1'b0,  10'd83},{ 8'd30, 1'b0, 10'd105},{ 8'd30, 1'b0, 10'd115},{ 8'd30, 1'b0, 10'd270},{ 8'd30, 1'b0, 10'd314},{ 8'd30, 1'b0, 10'd324},{ 8'd30, 1'b0, 10'd368},{ 8'd30, 1'b0, 10'd434},{ 8'd30, 1'b0, 10'd457},{ 8'd30, 1'b0, 10'd501},{ 8'd30, 1'b0, 10'd502},{ 8'd30, 1'b1, 10'd689},
{ 8'd29, 1'b0,  10'd61},{ 8'd29, 1'b0, 10'd159},{ 8'd29, 1'b0, 10'd181},{ 8'd29, 1'b0, 10'd193},{ 8'd29, 1'b0, 10'd247},{ 8'd29, 1'b0, 10'd335},{ 8'd29, 1'b0, 10'd435},{ 8'd29, 1'b0, 10'd468},{ 8'd29, 1'b0, 10'd556},{ 8'd29, 1'b0, 10'd611},{ 8'd29, 1'b0, 10'd690},{ 8'd29, 1'b1, 10'd731},
{ 8'd28, 1'b0,  10'd62},{ 8'd28, 1'b0, 10'd160},{ 8'd28, 1'b0, 10'd292},{ 8'd28, 1'b0, 10'd544},{ 8'd28, 1'b0, 10'd588},{ 8'd28, 1'b0, 10'd645},{ 8'd28, 1'b0, 10'd667},{ 8'd28, 1'b0, 10'd700},{ 8'd28, 1'b0, 10'd744},{ 8'd28, 1'b0, 10'd765},{ 8'd28, 1'b0, 10'd775},{ 8'd28, 1'b1, 10'd776},
{ 8'd27, 1'b0,  10'd38},{ 8'd27, 1'b0,  10'd84},{ 8'd27, 1'b0, 10'd172},{ 8'd27, 1'b0, 10'd182},{ 8'd27, 1'b0, 10'd215},{ 8'd27, 1'b0, 10'd258},{ 8'd27, 1'b0, 10'd259},{ 8'd27, 1'b0, 10'd260},{ 8'd27, 1'b0, 10'd325},{ 8'd27, 1'b0, 10'd390},{ 8'd27, 1'b0, 10'd533},{ 8'd27, 1'b1, 10'd612},
{ 8'd26, 1'b0,  10'd39},{ 8'd26, 1'b0, 10'd194},{ 8'd26, 1'b0, 10'd248},{ 8'd26, 1'b0, 10'd249},{ 8'd26, 1'b0, 10'd348},{ 8'd26, 1'b0, 10'd401},{ 8'd26, 1'b0, 10'd445},{ 8'd26, 1'b0, 10'd489},{ 8'd26, 1'b0, 10'd523},{ 8'd26, 1'b0, 10'd524},{ 8'd26, 1'b0, 10'd722},{ 8'd26, 1'b1, 10'd753},
{ 8'd25, 1'b0,  10'd49},{ 8'd25, 1'b0,  10'd63},{ 8'd25, 1'b0,  10'd71},{ 8'd25, 1'b0,  10'd85},{ 8'd25, 1'b0, 10'd139},{ 8'd25, 1'b0, 10'd281},{ 8'd25, 1'b0, 10'd425},{ 8'd25, 1'b0, 10'd446},{ 8'd25, 1'b0, 10'd458},{ 8'd25, 1'b0, 10'd459},{ 8'd25, 1'b0, 10'd646},{ 8'd25, 1'b1, 10'd668},
{ 8'd24, 1'b0,   10'd7},{ 8'd24, 1'b0,  10'd17},{ 8'd24, 1'b0,  10'd64},{ 8'd24, 1'b0, 10'd116},{ 8'd24, 1'b0, 10'd391},{ 8'd24, 1'b0, 10'd402},{ 8'd24, 1'b0, 10'd412},{ 8'd24, 1'b0, 10'd480},{ 8'd24, 1'b0, 10'd513},{ 8'd24, 1'b0, 10'd514},{ 8'd24, 1'b0, 10'd732},{ 8'd24, 1'b1, 10'd777},
{ 8'd23, 1'b0, 10'd117},{ 8'd23, 1'b0, 10'd173},{ 8'd23, 1'b0, 10'd195},{ 8'd23, 1'b0, 10'd203},{ 8'd23, 1'b0, 10'd226},{ 8'd23, 1'b0, 10'd358},{ 8'd23, 1'b0, 10'd379},{ 8'd23, 1'b0, 10'd380},{ 8'd23, 1'b0, 10'd545},{ 8'd23, 1'b0, 10'd568},{ 8'd23, 1'b0, 10'd578},{ 8'd23, 1'b1, 10'd711},
{ 8'd22, 1'b0,   10'd8},{ 8'd22, 1'b0,  10'd40},{ 8'd22, 1'b0,  10'd65},{ 8'd22, 1'b0,  10'd94},{ 8'd22, 1'b0, 10'd106},{ 8'd22, 1'b0, 10'd336},{ 8'd22, 1'b0, 10'd359},{ 8'd22, 1'b0, 10'd436},{ 8'd22, 1'b0, 10'd469},{ 8'd22, 1'b0, 10'd621},{ 8'd22, 1'b0, 10'd622},{ 8'd22, 1'b1, 10'd701},
{ 8'd21, 1'b0, 10'd250},{ 8'd21, 1'b0, 10'd271},{ 8'd21, 1'b0, 10'd360},{ 8'd21, 1'b0, 10'd525},{ 8'd21, 1'b0, 10'd534},{ 8'd21, 1'b0, 10'd535},{ 8'd21, 1'b0, 10'd579},{ 8'd21, 1'b0, 10'd580},{ 8'd21, 1'b0, 10'd676},{ 8'd21, 1'b0, 10'd733},{ 8'd21, 1'b0, 10'd787},{ 8'd21, 1'b1, 10'd788},
{ 8'd20, 1'b0,  10'd72},{ 8'd20, 1'b0, 10'd204},{ 8'd20, 1'b0, 10'd272},{ 8'd20, 1'b0, 10'd437},{ 8'd20, 1'b0, 10'd438},{ 8'd20, 1'b0, 10'd447},{ 8'd20, 1'b0, 10'd448},{ 8'd20, 1'b0, 10'd490},{ 8'd20, 1'b0, 10'd546},{ 8'd20, 1'b0, 10'd557},{ 8'd20, 1'b0, 10'd677},{ 8'd20, 1'b1, 10'd734},
{ 8'd19, 1'b0, 10'd183},{ 8'd19, 1'b0, 10'd227},{ 8'd19, 1'b0, 10'd261},{ 8'd19, 1'b0, 10'd381},{ 8'd19, 1'b0, 10'd413},{ 8'd19, 1'b0, 10'd600},{ 8'd19, 1'b0, 10'd633},{ 8'd19, 1'b0, 10'd654},{ 8'd19, 1'b0, 10'd735},{ 8'd19, 1'b0, 10'd766},{ 8'd19, 1'b0, 10'd778},{ 8'd19, 1'b1, 10'd789},
{ 8'd18, 1'b0,  10'd50},{ 8'd18, 1'b0,  10'd51},{ 8'd18, 1'b0,  10'd86},{ 8'd18, 1'b0, 10'd236},{ 8'd18, 1'b0, 10'd315},{ 8'd18, 1'b0, 10'd481},{ 8'd18, 1'b0, 10'd503},{ 8'd18, 1'b0, 10'd613},{ 8'd18, 1'b0, 10'd623},{ 8'd18, 1'b0, 10'd624},{ 8'd18, 1'b0, 10'd678},{ 8'd18, 1'b1, 10'd767},
{ 8'd17, 1'b0,  10'd41},{ 8'd17, 1'b0,  10'd42},{ 8'd17, 1'b0,  10'd73},{ 8'd17, 1'b0, 10'd118},{ 8'd17, 1'b0, 10'd161},{ 8'd17, 1'b0, 10'd251},{ 8'd17, 1'b0, 10'd282},{ 8'd17, 1'b0, 10'd293},{ 8'd17, 1'b0, 10'd414},{ 8'd17, 1'b0, 10'd601},{ 8'd17, 1'b0, 10'd723},{ 8'd17, 1'b1, 10'd754},
{ 8'd16, 1'b0, 10'd126},{ 8'd16, 1'b0, 10'd294},{ 8'd16, 1'b0, 10'd304},{ 8'd16, 1'b0, 10'd369},{ 8'd16, 1'b0, 10'd415},{ 8'd16, 1'b0, 10'd602},{ 8'd16, 1'b0, 10'd603},{ 8'd16, 1'b0, 10'd604},{ 8'd16, 1'b0, 10'd625},{ 8'd16, 1'b0, 10'd634},{ 8'd16, 1'b0, 10'd655},{ 8'd16, 1'b1, 10'd779},
{ 8'd15, 1'b0,   10'd9},{ 8'd15, 1'b0, 10'd127},{ 8'd15, 1'b0, 10'd150},{ 8'd15, 1'b0, 10'd162},{ 8'd15, 1'b0, 10'd174},{ 8'd15, 1'b0, 10'd184},{ 8'd15, 1'b0, 10'd237},{ 8'd15, 1'b0, 10'd439},{ 8'd15, 1'b0, 10'd449},{ 8'd15, 1'b0, 10'd491},{ 8'd15, 1'b0, 10'd626},{ 8'd15, 1'b1, 10'd790},
{ 8'd14, 1'b0,  10'd29},{ 8'd14, 1'b0,  10'd52},{ 8'd14, 1'b0, 10'd205},{ 8'd14, 1'b0, 10'd206},{ 8'd14, 1'b0, 10'd295},{ 8'd14, 1'b0, 10'd370},{ 8'd14, 1'b0, 10'd558},{ 8'd14, 1'b0, 10'd569},{ 8'd14, 1'b0, 10'd581},{ 8'd14, 1'b0, 10'd679},{ 8'd14, 1'b0, 10'd724},{ 8'd14, 1'b1, 10'd755},
{ 8'd13, 1'b0, 10'd119},{ 8'd13, 1'b0, 10'd140},{ 8'd13, 1'b0, 10'd163},{ 8'd13, 1'b0, 10'd185},{ 8'd13, 1'b0, 10'd337},{ 8'd13, 1'b0, 10'd392},{ 8'd13, 1'b0, 10'd403},{ 8'd13, 1'b0, 10'd526},{ 8'd13, 1'b0, 10'd536},{ 8'd13, 1'b0, 10'd547},{ 8'd13, 1'b0, 10'd589},{ 8'd13, 1'b1, 10'd780},
{ 8'd12, 1'b0,  10'd43},{ 8'd12, 1'b0,  10'd74},{ 8'd12, 1'b0, 10'd426},{ 8'd12, 1'b0, 10'd482},{ 8'd12, 1'b0, 10'd492},{ 8'd12, 1'b0, 10'd537},{ 8'd12, 1'b0, 10'd570},{ 8'd12, 1'b0, 10'd614},{ 8'd12, 1'b0, 10'd635},{ 8'd12, 1'b0, 10'd656},{ 8'd12, 1'b0, 10'd691},{ 8'd12, 1'b1, 10'd768},
{ 8'd11, 1'b0,  10'd18},{ 8'd11, 1'b0,  10'd53},{ 8'd11, 1'b0, 10'd107},{ 8'd11, 1'b0, 10'd128},{ 8'd11, 1'b0, 10'd129},{ 8'd11, 1'b0, 10'd141},{ 8'd11, 1'b0, 10'd228},{ 8'd11, 1'b0, 10'd283},{ 8'd11, 1'b0, 10'd326},{ 8'd11, 1'b0, 10'd427},{ 8'd11, 1'b0, 10'd450},{ 8'd11, 1'b1, 10'd769},
{ 8'd10, 1'b0,  10'd75},{ 8'd10, 1'b0,  10'd87},{ 8'd10, 1'b0, 10'd229},{ 8'd10, 1'b0, 10'd305},{ 8'd10, 1'b0, 10'd316},{ 8'd10, 1'b0, 10'd317},{ 8'd10, 1'b0, 10'd327},{ 8'd10, 1'b0, 10'd349},{ 8'd10, 1'b0, 10'd470},{ 8'd10, 1'b0, 10'd712},{ 8'd10, 1'b0, 10'd745},{ 8'd10, 1'b1, 10'd791},
{  8'd9, 1'b0,  10'd19},{  8'd9, 1'b0, 10'd130},{  8'd9, 1'b0, 10'd186},{  8'd9, 1'b0, 10'd216},{  8'd9, 1'b0, 10'd262},{  8'd9, 1'b0, 10'd428},{  8'd9, 1'b0, 10'd460},{  8'd9, 1'b0, 10'd504},{  8'd9, 1'b0, 10'd548},{  8'd9, 1'b0, 10'd590},{  8'd9, 1'b0, 10'd591},{  8'd9, 1'b1, 10'd636},
{  8'd8, 1'b0,  10'd30},{  8'd8, 1'b0,  10'd95},{  8'd8, 1'b0,  10'd96},{  8'd8, 1'b0,  10'd97},{  8'd8, 1'b0, 10'd338},{  8'd8, 1'b0, 10'd339},{  8'd8, 1'b0, 10'd371},{  8'd8, 1'b0, 10'd493},{  8'd8, 1'b0, 10'd494},{  8'd8, 1'b0, 10'd515},{  8'd8, 1'b0, 10'd516},{  8'd8, 1'b1, 10'd713},
{  8'd7, 1'b0,  10'd20},{  8'd7, 1'b0,  10'd54},{  8'd7, 1'b0, 10'd108},{  8'd7, 1'b0, 10'd151},{  8'd7, 1'b0, 10'd164},{  8'd7, 1'b0, 10'd217},{  8'd7, 1'b0, 10'd361},{  8'd7, 1'b0, 10'd527},{  8'd7, 1'b0, 10'd559},{  8'd7, 1'b0, 10'd582},{  8'd7, 1'b0, 10'd592},{  8'd7, 1'b1, 10'd725},
{  8'd6, 1'b0,  10'd31},{  8'd6, 1'b0,  10'd76},{  8'd6, 1'b0, 10'd238},{  8'd6, 1'b0, 10'd273},{  8'd6, 1'b0, 10'd306},{  8'd6, 1'b0, 10'd362},{  8'd6, 1'b0, 10'd382},{  8'd6, 1'b0, 10'd669},{  8'd6, 1'b0, 10'd714},{  8'd6, 1'b0, 10'd746},{  8'd6, 1'b0, 10'd747},{  8'd6, 1'b1, 10'd756},
{  8'd5, 1'b0, 10'd142},{  8'd5, 1'b0, 10'd196},{  8'd5, 1'b0, 10'd218},{  8'd5, 1'b0, 10'd328},{  8'd5, 1'b0, 10'd404},{  8'd5, 1'b0, 10'd416},{  8'd5, 1'b0, 10'd560},{  8'd5, 1'b0, 10'd647},{  8'd5, 1'b0, 10'd657},{  8'd5, 1'b0, 10'd680},{  8'd5, 1'b0, 10'd736},{  8'd5, 1'b1, 10'd757},
{  8'd4, 1'b0, 10'd131},{  8'd4, 1'b0, 10'd175},{  8'd4, 1'b0, 10'd207},{  8'd4, 1'b0, 10'd239},{  8'd4, 1'b0, 10'd350},{  8'd4, 1'b0, 10'd405},{  8'd4, 1'b0, 10'd461},{  8'd4, 1'b0, 10'd483},{  8'd4, 1'b0, 10'd538},{  8'd4, 1'b0, 10'd658},{  8'd4, 1'b0, 10'd702},{  8'd4, 1'b1, 10'd758},
{  8'd3, 1'b0,  10'd98},{  8'd3, 1'b0, 10'd152},{  8'd3, 1'b0, 10'd153},{  8'd3, 1'b0, 10'd240},{  8'd3, 1'b0, 10'd252},{  8'd3, 1'b0, 10'd372},{  8'd3, 1'b0, 10'd383},{  8'd3, 1'b0, 10'd393},{  8'd3, 1'b0, 10'd394},{  8'd3, 1'b0, 10'd549},{  8'd3, 1'b0, 10'd659},{  8'd3, 1'b1, 10'd681},
{  8'd2, 1'b0,  10'd32},{  8'd2, 1'b0, 10'd197},{  8'd2, 1'b0, 10'd219},{  8'd2, 1'b0, 10'd230},{  8'd2, 1'b0, 10'd241},{  8'd2, 1'b0, 10'd318},{  8'd2, 1'b0, 10'd329},{  8'd2, 1'b0, 10'd373},{  8'd2, 1'b0, 10'd471},{  8'd2, 1'b0, 10'd505},{  8'd2, 1'b0, 10'd637},{  8'd2, 1'b1, 10'd670},
{  8'd1, 1'b0, 10'd120},{  8'd1, 1'b0, 10'd208},{  8'd1, 1'b0, 10'd263},{  8'd1, 1'b0, 10'd274},{  8'd1, 1'b0, 10'd284},{  8'd1, 1'b0, 10'd285},{  8'd1, 1'b0, 10'd351},{  8'd1, 1'b0, 10'd406},{  8'd1, 1'b0, 10'd417},{  8'd1, 1'b0, 10'd571},{  8'd1, 1'b0, 10'd615},{  8'd1, 1'b1, 10'd703},
{  8'd0, 1'b0,  10'd10},{  8'd0, 1'b0,  10'd21},{  8'd0, 1'b0, 10'd109},{  8'd0, 1'b0, 10'd296},{  8'd0, 1'b0, 10'd307},{  8'd0, 1'b0, 10'd340},{  8'd0, 1'b0, 10'd384},{  8'd0, 1'b0, 10'd395},{  8'd0, 1'b0, 10'd472},{  8'd0, 1'b0, 10'd593},{  8'd0, 1'b0, 10'd648},{  8'd0, 1'b1, 10'd692}
};
localparam int          cLARGE_HS_TAB_2BY3_PACKED_SIZE = 600;
localparam bit [18 : 0] cLARGE_HS_TAB_2BY3_PACKED[cLARGE_HS_TAB_2BY3_PACKED_SIZE] = '{
{  1'b1, 1'b0, 8'd179,    9'd1},{  1'b0, 1'b0, 8'd120,    9'd0},{  1'b0, 1'b0,  8'd79,  9'd232},{  1'b0, 1'b0,  8'd79,  9'd165},{  1'b0, 1'b0,  8'd60,    9'd0},{  1'b0, 1'b0,  8'd39,  9'd284},{  1'b0, 1'b0,  8'd12,  9'd230},{  1'b0, 1'b0,  8'd11,  9'd236},{  1'b0, 1'b0,   8'd0,    9'd0},{  1'b0, 1'b1,   8'd0,    9'd4},
{  1'b0, 1'b0, 8'd121,    9'd0},{  1'b0, 1'b0, 8'd120,    9'd0},{  1'b0, 1'b0, 8'd112,  9'd302},{  1'b0, 1'b0, 8'd111,   9'd61},{  1'b0, 1'b0,  8'd61,    9'd0},{  1'b0, 1'b0,  8'd17,  9'd225},{  1'b0, 1'b0,  8'd12,  9'd236},{  1'b0, 1'b0,   8'd7,  9'd311},{  1'b0, 1'b0,   8'd3,  9'd189},{  1'b0, 1'b1,   8'd1,    9'd0},
{  1'b0, 1'b0, 8'd122,    9'd0},{  1'b0, 1'b0, 8'd121,    9'd0},{  1'b0, 1'b0, 8'd117,  9'd112},{  1'b0, 1'b0,  8'd85,   9'd72},{  1'b0, 1'b0,  8'd62,    9'd0},{  1'b0, 1'b0,  8'd47,  9'd351},{  1'b0, 1'b0,  8'd39,  9'd318},{  1'b0, 1'b0,  8'd11,   9'd72},{  1'b0, 1'b0,   8'd8,  9'd151},{  1'b0, 1'b1,   8'd2,    9'd0},
{  1'b0, 1'b0, 8'd123,    9'd0},{  1'b0, 1'b0, 8'd122,    9'd0},{  1'b0, 1'b0, 8'd114,  9'd300},{  1'b0, 1'b0, 8'd106,  9'd267},{  1'b0, 1'b0,  8'd63,    9'd0},{  1'b0, 1'b0,  8'd16,   9'd19},{  1'b0, 1'b0,   8'd6,  9'd229},{  1'b0, 1'b0,   8'd3,    9'd0},{  1'b0, 1'b0,   8'd3,  9'd103},{  1'b0, 1'b1,   8'd1,  9'd308},
{  1'b0, 1'b0, 8'd124,    9'd0},{  1'b0, 1'b0, 8'd123,    9'd0},{  1'b0, 1'b0,  8'd78,   9'd34},{  1'b0, 1'b0,  8'd72,  9'd266},{  1'b0, 1'b0,  8'd64,    9'd0},{  1'b0, 1'b0,  8'd58,   9'd31},{  1'b0, 1'b0,  8'd30,  9'd339},{  1'b0, 1'b0,   8'd4,    9'd0},{  1'b0, 1'b0,   8'd2,  9'd201},{  1'b0, 1'b1,   8'd1,   9'd97},
{  1'b0, 1'b0, 8'd125,    9'd0},{  1'b0, 1'b0, 8'd124,    9'd0},{  1'b0, 1'b0,  8'd66,  9'd193},{  1'b0, 1'b0,  8'd65,    9'd0},{  1'b0, 1'b0,  8'd62,   9'd51},{  1'b0, 1'b0,  8'd57,  9'd164},{  1'b0, 1'b0,   8'd9,  9'd158},{  1'b0, 1'b0,   8'd7,   9'd92},{  1'b0, 1'b0,   8'd5,    9'd0},{  1'b0, 1'b1,   8'd5,  9'd312},
{  1'b0, 1'b0, 8'd126,    9'd0},{  1'b0, 1'b0, 8'd125,    9'd0},{  1'b0, 1'b0,  8'd83,  9'd162},{  1'b0, 1'b0,  8'd69,   9'd20},{  1'b0, 1'b0,  8'd66,    9'd0},{  1'b0, 1'b0,  8'd35,   9'd96},{  1'b0, 1'b0,   8'd8,  9'd213},{  1'b0, 1'b0,   8'd6,    9'd0},{  1'b0, 1'b0,   8'd6,    9'd8},{  1'b0, 1'b1,   8'd0,  9'd137},
{  1'b0, 1'b0, 8'd127,    9'd0},{  1'b0, 1'b0, 8'd126,    9'd0},{  1'b0, 1'b0,  8'd99,  9'd286},{  1'b0, 1'b0,  8'd88,  9'd123},{  1'b0, 1'b0,  8'd67,    9'd0},{  1'b0, 1'b0,  8'd14,  9'd267},{  1'b0, 1'b0,   8'd7,    9'd0},{  1'b0, 1'b0,   8'd7,  9'd344},{  1'b0, 1'b0,   8'd1,  9'd224},{  1'b0, 1'b1,   8'd0,   9'd46},
{  1'b0, 1'b0, 8'd128,    9'd0},{  1'b0, 1'b0, 8'd127,    9'd0},{  1'b0, 1'b0, 8'd110,  9'd269},{  1'b0, 1'b0, 8'd107,   9'd84},{  1'b0, 1'b0,  8'd68,    9'd0},{  1'b0, 1'b0,  8'd31,  9'd243},{  1'b0, 1'b0,  8'd13,   9'd49},{  1'b0, 1'b0,  8'd11,  9'd210},{  1'b0, 1'b0,  8'd10,    9'd6},{  1'b0, 1'b1,   8'd8,    9'd0},
{  1'b0, 1'b0, 8'd129,    9'd0},{  1'b0, 1'b0, 8'd128,    9'd0},{  1'b0, 1'b0, 8'd103,  9'd307},{  1'b0, 1'b0,  8'd94,   9'd26},{  1'b0, 1'b0,  8'd69,    9'd0},{  1'b0, 1'b0,  8'd42,  9'd104},{  1'b0, 1'b0,   8'd9,    9'd0},{  1'b0, 1'b0,   8'd7,  9'd176},{  1'b0, 1'b0,   8'd5,  9'd206},{  1'b0, 1'b1,   8'd4,  9'd328},
{  1'b0, 1'b0, 8'd130,    9'd0},{  1'b0, 1'b0, 8'd129,    9'd0},{  1'b0, 1'b0,  8'd94,  9'd125},{  1'b0, 1'b0,  8'd85,  9'd133},{  1'b0, 1'b0,  8'd70,    9'd0},{  1'b0, 1'b0,  8'd42,  9'd317},{  1'b0, 1'b0,  8'd38,   9'd68},{  1'b0, 1'b0,  8'd10,    9'd0},{  1'b0, 1'b0,   8'd7,  9'd135},{  1'b0, 1'b1,   8'd6,  9'd207},
{  1'b0, 1'b0, 8'd131,    9'd0},{  1'b0, 1'b0, 8'd130,    9'd0},{  1'b0, 1'b0,  8'd97,    9'd3},{  1'b0, 1'b0,  8'd82,  9'd102},{  1'b0, 1'b0,  8'd71,    9'd0},{  1'b0, 1'b0,  8'd33,  9'd324},{  1'b0, 1'b0,  8'd11,    9'd0},{  1'b0, 1'b0,   8'd8,   9'd63},{  1'b0, 1'b0,   8'd6,   9'd93},{  1'b0, 1'b1,   8'd2,  9'd119},
{  1'b0, 1'b0, 8'd132,    9'd0},{  1'b0, 1'b0, 8'd131,    9'd0},{  1'b0, 1'b0, 8'd103,  9'd141},{  1'b0, 1'b0,  8'd72,    9'd0},{  1'b0, 1'b0,  8'd63,  9'd304},{  1'b0, 1'b0,  8'd56,   9'd40},{  1'b0, 1'b0,  8'd44,  9'd196},{  1'b0, 1'b0,  8'd12,    9'd0},{  1'b0, 1'b0,   8'd9,  9'd337},{  1'b0, 1'b1,   8'd3,  9'd166},
{  1'b0, 1'b0, 8'd133,    9'd0},{  1'b0, 1'b0, 8'd132,    9'd0},{  1'b0, 1'b0,  8'd76,    9'd4},{  1'b0, 1'b0,  8'd73,    9'd0},{  1'b0, 1'b0,  8'd65,  9'd169},{  1'b0, 1'b0,  8'd40,  9'd337},{  1'b0, 1'b0,  8'd13,    9'd0},{  1'b0, 1'b0,  8'd11,   9'd67},{  1'b0, 1'b0,   8'd1,  9'd107},{  1'b0, 1'b1,   8'd0,  9'd311},
{  1'b0, 1'b0, 8'd134,    9'd0},{  1'b0, 1'b0, 8'd133,    9'd0},{  1'b0, 1'b0,  8'd82,   9'd90},{  1'b0, 1'b0,  8'd77,   9'd21},{  1'b0, 1'b0,  8'd74,    9'd0},{  1'b0, 1'b0,  8'd27,  9'd273},{  1'b0, 1'b0,  8'd23,  9'd210},{  1'b0, 1'b0,  8'd14,    9'd0},{  1'b0, 1'b0,   8'd4,  9'd298},{  1'b0, 1'b1,   8'd2,  9'd213},
{  1'b0, 1'b0, 8'd135,    9'd0},{  1'b0, 1'b0, 8'd134,    9'd0},{  1'b0, 1'b0, 8'd107,  9'd293},{  1'b0, 1'b0,  8'd75,    9'd0},{  1'b0, 1'b0,  8'd71,  9'd156},{  1'b0, 1'b0,  8'd56,  9'd288},{  1'b0, 1'b0,  8'd25,  9'd293},{  1'b0, 1'b0,  8'd15,    9'd0},{  1'b0, 1'b0,  8'd10,   9'd15},{  1'b0, 1'b1,   8'd2,   9'd74},
{  1'b0, 1'b0, 8'd136,    9'd0},{  1'b0, 1'b0, 8'd135,    9'd0},{  1'b0, 1'b0, 8'd102,   9'd84},{  1'b0, 1'b0,  8'd86,  9'd260},{  1'b0, 1'b0,  8'd76,    9'd0},{  1'b0, 1'b0,  8'd34,    9'd8},{  1'b0, 1'b0,  8'd19,  9'd359},{  1'b0, 1'b0,  8'd16,    9'd0},{  1'b0, 1'b0,  8'd10,  9'd226},{  1'b0, 1'b1,   8'd3,  9'd242},
{  1'b0, 1'b0, 8'd137,    9'd0},{  1'b0, 1'b0, 8'd136,    9'd0},{  1'b0, 1'b0, 8'd108,   9'd80},{  1'b0, 1'b0,  8'd78,  9'd246},{  1'b0, 1'b0,  8'd77,    9'd0},{  1'b0, 1'b0,  8'd34,   9'd70},{  1'b0, 1'b0,  8'd17,    9'd0},{  1'b0, 1'b0,   8'd6,  9'd192},{  1'b0, 1'b0,   8'd5,   9'd33},{  1'b0, 1'b1,   8'd2,  9'd299},
{  1'b0, 1'b0, 8'd138,    9'd0},{  1'b0, 1'b0, 8'd137,    9'd0},{  1'b0, 1'b0,  8'd88,  9'd345},{  1'b0, 1'b0,  8'd78,    9'd0},{  1'b0, 1'b0,  8'd66,  9'd151},{  1'b0, 1'b0,  8'd38,   9'd97},{  1'b0, 1'b0,  8'd29,  9'd111},{  1'b0, 1'b0,  8'd18,    9'd0},{  1'b0, 1'b0,   8'd9,  9'd275},{  1'b0, 1'b1,   8'd5,  9'd253},
{  1'b0, 1'b0, 8'd139,    9'd0},{  1'b0, 1'b0, 8'd138,    9'd0},{  1'b0, 1'b0,  8'd84,   9'd91},{  1'b0, 1'b0,  8'd79,    9'd0},{  1'b0, 1'b0,  8'd67,   9'd89},{  1'b0, 1'b0,  8'd50,   9'd55},{  1'b0, 1'b0,  8'd47,  9'd196},{  1'b0, 1'b0,  8'd19,    9'd0},{  1'b0, 1'b0,   8'd9,  9'd333},{  1'b0, 1'b1,   8'd0,  9'd176},
{  1'b0, 1'b0, 8'd140,    9'd0},{  1'b0, 1'b0, 8'd139,    9'd0},{  1'b0, 1'b0,  8'd90,   9'd43},{  1'b0, 1'b0,  8'd80,    9'd0},{  1'b0, 1'b0,  8'd61,  9'd156},{  1'b0, 1'b0,  8'd44,  9'd329},{  1'b0, 1'b0,  8'd20,    9'd0},{  1'b0, 1'b0,  8'd16,  9'd150},{  1'b0, 1'b0,   8'd5,   9'd28},{  1'b0, 1'b1,   8'd1,   9'd85},
{  1'b0, 1'b0, 8'd141,    9'd0},{  1'b0, 1'b0, 8'd140,    9'd0},{  1'b0, 1'b0,  8'd87,  9'd259},{  1'b0, 1'b0,  8'd81,    9'd0},{  1'b0, 1'b0,  8'd81,  9'd165},{  1'b0, 1'b0,  8'd36,  9'd175},{  1'b0, 1'b0,  8'd28,  9'd116},{  1'b0, 1'b0,  8'd21,    9'd0},{  1'b0, 1'b0,   8'd7,  9'd202},{  1'b0, 1'b1,   8'd7,  9'd307},
{  1'b0, 1'b0, 8'd142,    9'd0},{  1'b0, 1'b0, 8'd141,    9'd0},{  1'b0, 1'b0,  8'd82,    9'd0},{  1'b0, 1'b0,  8'd74,  9'd133},{  1'b0, 1'b0,  8'd70,   9'd18},{  1'b0, 1'b0,  8'd55,   9'd86},{  1'b0, 1'b0,  8'd48,  9'd161},{  1'b0, 1'b0,  8'd22,    9'd0},{  1'b0, 1'b0,   8'd8,  9'd161},{  1'b0, 1'b1,   8'd3,  9'd136},
{  1'b0, 1'b0, 8'd143,    9'd0},{  1'b0, 1'b0, 8'd142,    9'd0},{  1'b0, 1'b0, 8'd115,   9'd88},{  1'b0, 1'b0, 8'd115,   9'd51},{  1'b0, 1'b0,  8'd83,    9'd0},{  1'b0, 1'b0,  8'd53,   9'd99},{  1'b0, 1'b0,  8'd23,    9'd0},{  1'b0, 1'b0,  8'd11,  9'd170},{  1'b0, 1'b0,   8'd4,  9'd102},{  1'b0, 1'b1,   8'd0,  9'd267},
{  1'b0, 1'b0, 8'd144,    9'd0},{  1'b0, 1'b0, 8'd143,    9'd0},{  1'b0, 1'b0,  8'd89,  9'd313},{  1'b0, 1'b0,  8'd84,    9'd0},{  1'b0, 1'b0,  8'd68,  9'd150},{  1'b0, 1'b0,  8'd45,  9'd327},{  1'b0, 1'b0,  8'd24,    9'd0},{  1'b0, 1'b0,  8'd11,  9'd358},{  1'b0, 1'b0,   8'd8,  9'd254},{  1'b0, 1'b1,   8'd2,  9'd100},
{  1'b0, 1'b0, 8'd145,    9'd0},{  1'b0, 1'b0, 8'd144,    9'd0},{  1'b0, 1'b0, 8'd105,  9'd272},{  1'b0, 1'b0,  8'd98,  9'd311},{  1'b0, 1'b0,  8'd85,    9'd0},{  1'b0, 1'b0,  8'd37,  9'd198},{  1'b0, 1'b0,  8'd25,    9'd0},{  1'b0, 1'b0,   8'd9,  9'd325},{  1'b0, 1'b0,   8'd1,  9'd230},{  1'b0, 1'b1,   8'd0,  9'd134},
{  1'b0, 1'b0, 8'd146,    9'd0},{  1'b0, 1'b0, 8'd145,    9'd0},{  1'b0, 1'b0,  8'd86,    9'd0},{  1'b0, 1'b0,  8'd81,  9'd303},{  1'b0, 1'b0,  8'd77,  9'd321},{  1'b0, 1'b0,  8'd54,  9'd122},{  1'b0, 1'b0,  8'd54,  9'd195},{  1'b0, 1'b0,  8'd26,    9'd0},{  1'b0, 1'b0,   8'd4,   9'd88},{  1'b0, 1'b1,   8'd0,    9'd8},
{  1'b0, 1'b0, 8'd147,    9'd0},{  1'b0, 1'b0, 8'd146,    9'd0},{  1'b0, 1'b0,  8'd96,  9'd152},{  1'b0, 1'b0,  8'd87,    9'd0},{  1'b0, 1'b0,  8'd72,  9'd100},{  1'b0, 1'b0,  8'd58,  9'd111},{  1'b0, 1'b0,  8'd30,  9'd216},{  1'b0, 1'b0,  8'd27,    9'd0},{  1'b0, 1'b0,   8'd4,  9'd278},{  1'b0, 1'b1,   8'd1,  9'd286},
{  1'b0, 1'b0, 8'd148,    9'd0},{  1'b0, 1'b0, 8'd147,    9'd0},{  1'b0, 1'b0, 8'd113,  9'd149},{  1'b0, 1'b0, 8'd105,  9'd212},{  1'b0, 1'b0,  8'd88,    9'd0},{  1'b0, 1'b0,  8'd28,    9'd0},{  1'b0, 1'b0,  8'd22,  9'd167},{  1'b0, 1'b0,  8'd10,   9'd76},{  1'b0, 1'b0,  8'd10,   9'd58},{  1'b0, 1'b1,   8'd2,  9'd310},
{  1'b0, 1'b0, 8'd149,    9'd0},{  1'b0, 1'b0, 8'd148,    9'd0},{  1'b0, 1'b0,  8'd91,  9'd298},{  1'b0, 1'b0,  8'd89,    9'd0},{  1'b0, 1'b0,  8'd73,  9'd246},{  1'b0, 1'b0,  8'd55,   9'd93},{  1'b0, 1'b0,  8'd29,    9'd0},{  1'b0, 1'b0,  8'd28,  9'd123},{  1'b0, 1'b0,  8'd11,  9'd137},{  1'b0, 1'b1,   8'd9,  9'd153},
{  1'b0, 1'b0, 8'd150,    9'd0},{  1'b0, 1'b0, 8'd149,    9'd0},{  1'b0, 1'b0,  8'd97,  9'd277},{  1'b0, 1'b0,  8'd90,    9'd0},{  1'b0, 1'b0,  8'd86,   9'd92},{  1'b0, 1'b0,  8'd35,  9'd121},{  1'b0, 1'b0,  8'd30,    9'd0},{  1'b0, 1'b0,  8'd18,   9'd36},{  1'b0, 1'b0,   8'd9,  9'd111},{  1'b0, 1'b1,   8'd5,  9'd281},
{  1'b0, 1'b0, 8'd151,    9'd0},{  1'b0, 1'b0, 8'd150,    9'd0},{  1'b0, 1'b0, 8'd117,   9'd79},{  1'b0, 1'b0, 8'd100,   9'd56},{  1'b0, 1'b0,  8'd91,    9'd0},{  1'b0, 1'b0,  8'd31,    9'd0},{  1'b0, 1'b0,  8'd11,   9'd10},{  1'b0, 1'b0,   8'd7,  9'd238},{  1'b0, 1'b0,   8'd6,  9'd290},{  1'b0, 1'b1,   8'd4,   9'd77},
{  1'b0, 1'b0, 8'd152,    9'd0},{  1'b0, 1'b0, 8'd151,    9'd0},{  1'b0, 1'b0,  8'd92,    9'd0},{  1'b0, 1'b0,  8'd80,    9'd7},{  1'b0, 1'b0,  8'd73,  9'd107},{  1'b0, 1'b0,  8'd32,    9'd0},{  1'b0, 1'b0,  8'd11,  9'd234},{  1'b0, 1'b0,   8'd7,  9'd136},{  1'b0, 1'b0,   8'd5,   9'd42},{  1'b0, 1'b1,   8'd1,  9'd213},
{  1'b0, 1'b0, 8'd153,    9'd0},{  1'b0, 1'b0, 8'd152,    9'd0},{  1'b0, 1'b0, 8'd113,  9'd196},{  1'b0, 1'b0, 8'd104,  9'd201},{  1'b0, 1'b0,  8'd93,    9'd0},{  1'b0, 1'b0,  8'd33,    9'd0},{  1'b0, 1'b0,  8'd26,   9'd98},{  1'b0, 1'b0,  8'd10,  9'd184},{  1'b0, 1'b0,   8'd9,  9'd122},{  1'b0, 1'b1,   8'd1,  9'd138},
{  1'b0, 1'b0, 8'd154,    9'd0},{  1'b0, 1'b0, 8'd153,    9'd0},{  1'b0, 1'b0,  8'd94,    9'd0},{  1'b0, 1'b0,  8'd69,  9'd272},{  1'b0, 1'b0,  8'd65,  9'd178},{  1'b0, 1'b0,  8'd57,  9'd341},{  1'b0, 1'b0,  8'd52,  9'd131},{  1'b0, 1'b0,  8'd34,    9'd0},{  1'b0, 1'b0,   8'd7,  9'd195},{  1'b0, 1'b1,   8'd3,  9'd290},
{  1'b0, 1'b0, 8'd155,    9'd0},{  1'b0, 1'b0, 8'd154,    9'd0},{  1'b0, 1'b0, 8'd108,  9'd316},{  1'b0, 1'b0,  8'd95,    9'd0},{  1'b0, 1'b0,  8'd68,  9'd158},{  1'b0, 1'b0,  8'd35,    9'd0},{  1'b0, 1'b0,  8'd26,  9'd141},{  1'b0, 1'b0,  8'd23,    9'd8},{  1'b0, 1'b0,  8'd11,  9'd206},{  1'b0, 1'b1,   8'd2,   9'd98},
{  1'b0, 1'b0, 8'd156,    9'd0},{  1'b0, 1'b0, 8'd155,    9'd0},{  1'b0, 1'b0,  8'd96,    9'd0},{  1'b0, 1'b0,  8'd91,  9'd108},{  1'b0, 1'b0,  8'd71,  9'd346},{  1'b0, 1'b0,  8'd51,   9'd72},{  1'b0, 1'b0,  8'd36,    9'd0},{  1'b0, 1'b0,  8'd19,  9'd203},{  1'b0, 1'b0,   8'd5,  9'd201},{  1'b0, 1'b1,   8'd3,   9'd92},
{  1'b0, 1'b0, 8'd157,    9'd0},{  1'b0, 1'b0, 8'd156,    9'd0},{  1'b0, 1'b0,  8'd99,  9'd348},{  1'b0, 1'b0,  8'd98,  9'd259},{  1'b0, 1'b0,  8'd97,    9'd0},{  1'b0, 1'b0,  8'd37,    9'd0},{  1'b0, 1'b0,  8'd20,  9'd331},{  1'b0, 1'b0,   8'd9,  9'd129},{  1'b0, 1'b0,   8'd3,  9'd329},{  1'b0, 1'b1,   8'd2,  9'd340},
{  1'b0, 1'b0, 8'd158,    9'd0},{  1'b0, 1'b0, 8'd157,    9'd0},{  1'b0, 1'b0, 8'd102,  9'd153},{  1'b0, 1'b0,  8'd98,    9'd0},{  1'b0, 1'b0,  8'd92,    9'd1},{  1'b0, 1'b0,  8'd38,    9'd0},{  1'b0, 1'b0,  8'd32,  9'd298},{  1'b0, 1'b0,  8'd21,  9'd132},{  1'b0, 1'b0,   8'd9,  9'd139},{  1'b0, 1'b1,   8'd4,  9'd243},
{  1'b0, 1'b0, 8'd159,    9'd0},{  1'b0, 1'b0, 8'd158,    9'd0},{  1'b0, 1'b0, 8'd111,   9'd50},{  1'b0, 1'b0,  8'd99,    9'd0},{  1'b0, 1'b0,  8'd93,  9'd342},{  1'b0, 1'b0,  8'd39,    9'd0},{  1'b0, 1'b0,  8'd37,  9'd339},{  1'b0, 1'b0,  8'd29,  9'd265},{  1'b0, 1'b0,  8'd11,  9'd332},{  1'b0, 1'b1,   8'd0,  9'd154},
{  1'b0, 1'b0, 8'd160,    9'd0},{  1'b0, 1'b0, 8'd159,    9'd0},{  1'b0, 1'b0, 8'd118,  9'd132},{  1'b0, 1'b0, 8'd100,    9'd0},{  1'b0, 1'b0,  8'd95,  9'd266},{  1'b0, 1'b0,  8'd53,   9'd72},{  1'b0, 1'b0,  8'd40,    9'd0},{  1'b0, 1'b0,  8'd22,  9'd265},{  1'b0, 1'b0,   8'd7,   9'd69},{  1'b0, 1'b1,   8'd1,  9'd165},
{  1'b0, 1'b0, 8'd161,    9'd0},{  1'b0, 1'b0, 8'd160,    9'd0},{  1'b0, 1'b0, 8'd101,    9'd0},{  1'b0, 1'b0,  8'd87,  9'd177},{  1'b0, 1'b0,  8'd64,  9'd152},{  1'b0, 1'b0,  8'd46,   9'd58},{  1'b0, 1'b0,  8'd41,    9'd0},{  1'b0, 1'b0,  8'd24,  9'd141},{  1'b0, 1'b0,   8'd7,  9'd262},{  1'b0, 1'b1,   8'd2,  9'd144},
{  1'b0, 1'b0, 8'd162,    9'd0},{  1'b0, 1'b0, 8'd161,    9'd0},{  1'b0, 1'b0, 8'd102,    9'd0},{  1'b0, 1'b0,  8'd75,  9'd245},{  1'b0, 1'b0,  8'd64,  9'd260},{  1'b0, 1'b0,  8'd48,  9'd217},{  1'b0, 1'b0,  8'd42,    9'd0},{  1'b0, 1'b0,  8'd15,  9'd184},{  1'b0, 1'b0,  8'd10,  9'd336},{  1'b0, 1'b1,   8'd5,  9'd264},
{  1'b0, 1'b0, 8'd163,    9'd0},{  1'b0, 1'b0, 8'd162,    9'd0},{  1'b0, 1'b0, 8'd109,  9'd274},{  1'b0, 1'b0, 8'd103,    9'd0},{  1'b0, 1'b0,  8'd96,  9'd171},{  1'b0, 1'b0,  8'd43,    9'd0},{  1'b0, 1'b0,  8'd33,  9'd111},{  1'b0, 1'b0,  8'd27,  9'd173},{  1'b0, 1'b0,   8'd9,   9'd52},{  1'b0, 1'b1,   8'd6,   9'd24},
{  1'b0, 1'b0, 8'd164,    9'd0},{  1'b0, 1'b0, 8'd163,    9'd0},{  1'b0, 1'b0, 8'd104,    9'd0},{  1'b0, 1'b0,  8'd93,   9'd61},{  1'b0, 1'b0,  8'd90,  9'd149},{  1'b0, 1'b0,  8'd59,  9'd342},{  1'b0, 1'b0,  8'd44,    9'd0},{  1'b0, 1'b0,  8'd25,  9'd279},{  1'b0, 1'b0,   8'd4,  9'd344},{  1'b0, 1'b1,   8'd1,  9'd103},
{  1'b0, 1'b0, 8'd165,    9'd0},{  1'b0, 1'b0, 8'd164,    9'd0},{  1'b0, 1'b0, 8'd105,    9'd0},{  1'b0, 1'b0,  8'd84,  9'd200},{  1'b0, 1'b0,  8'd76,   9'd50},{  1'b0, 1'b0,  8'd45,    9'd0},{  1'b0, 1'b0,  8'd41,  9'd322},{  1'b0, 1'b0,  8'd36,  9'd148},{  1'b0, 1'b0,  8'd10,  9'd181},{  1'b0, 1'b1,   8'd6,  9'd235},
{  1'b0, 1'b0, 8'd166,    9'd0},{  1'b0, 1'b0, 8'd165,    9'd0},{  1'b0, 1'b0, 8'd106,    9'd0},{  1'b0, 1'b0,  8'd61,  9'd137},{  1'b0, 1'b0,  8'd60,  9'd303},{  1'b0, 1'b0,  8'd46,    9'd0},{  1'b0, 1'b0,  8'd41,  9'd325},{  1'b0, 1'b0,  8'd15,  9'd341},{  1'b0, 1'b0,   8'd8,  9'd320},{  1'b0, 1'b1,   8'd0,  9'd213},
{  1'b0, 1'b0, 8'd167,    9'd0},{  1'b0, 1'b0, 8'd166,    9'd0},{  1'b0, 1'b0, 8'd114,  9'd223},{  1'b0, 1'b0, 8'd107,    9'd0},{  1'b0, 1'b0,  8'd60,  9'd286},{  1'b0, 1'b0,  8'd50,  9'd184},{  1'b0, 1'b0,  8'd47,    9'd0},{  1'b0, 1'b0,  8'd13,  9'd160},{  1'b0, 1'b0,   8'd6,  9'd253},{  1'b0, 1'b1,   8'd6,   9'd64},
{  1'b0, 1'b0, 8'd168,    9'd0},{  1'b0, 1'b0, 8'd167,    9'd0},{  1'b0, 1'b0, 8'd116,  9'd277},{  1'b0, 1'b0, 8'd108,    9'd0},{  1'b0, 1'b0,  8'd92,  9'd185},{  1'b0, 1'b0,  8'd48,    9'd0},{  1'b0, 1'b0,  8'd45,  9'd123},{  1'b0, 1'b0,  8'd18,   9'd25},{  1'b0, 1'b0,   8'd4,   9'd26},{  1'b0, 1'b1,   8'd0,  9'd348},
{  1'b0, 1'b0, 8'd169,    9'd0},{  1'b0, 1'b0, 8'd168,    9'd0},{  1'b0, 1'b0, 8'd119,   9'd59},{  1'b0, 1'b0, 8'd109,    9'd0},{  1'b0, 1'b0,  8'd75,  9'd234},{  1'b0, 1'b0,  8'd49,    9'd0},{  1'b0, 1'b0,  8'd21,   9'd69},{  1'b0, 1'b0,  8'd10,  9'd111},{  1'b0, 1'b0,   8'd5,   9'd51},{  1'b0, 1'b1,   8'd3,  9'd295},
{  1'b0, 1'b0, 8'd170,    9'd0},{  1'b0, 1'b0, 8'd169,    9'd0},{  1'b0, 1'b0, 8'd119,  9'd243},{  1'b0, 1'b0, 8'd112,  9'd316},{  1'b0, 1'b0, 8'd110,    9'd0},{  1'b0, 1'b0,  8'd50,    9'd0},{  1'b0, 1'b0,  8'd31,   9'd41},{  1'b0, 1'b0,  8'd24,  9'd140},{  1'b0, 1'b0,   8'd8,  9'd166},{  1'b0, 1'b1,   8'd2,  9'd182},
{  1'b0, 1'b0, 8'd171,    9'd0},{  1'b0, 1'b0, 8'd170,    9'd0},{  1'b0, 1'b0, 8'd116,    9'd8},{  1'b0, 1'b0, 8'd111,    9'd0},{  1'b0, 1'b0,  8'd74,  9'd309},{  1'b0, 1'b0,  8'd51,    9'd0},{  1'b0, 1'b0,  8'd10,  9'd352},{  1'b0, 1'b0,   8'd6,  9'd101},{  1'b0, 1'b0,   8'd5,   9'd80},{  1'b0, 1'b1,   8'd0,  9'd174},
{  1'b0, 1'b0, 8'd172,    9'd0},{  1'b0, 1'b0, 8'd171,    9'd0},{  1'b0, 1'b0, 8'd112,    9'd0},{  1'b0, 1'b0, 8'd101,  9'd334},{  1'b0, 1'b0,  8'd95,  9'd194},{  1'b0, 1'b0,  8'd52,    9'd0},{  1'b0, 1'b0,  8'd51,  9'd314},{  1'b0, 1'b0,  8'd40,  9'd205},{  1'b0, 1'b0,   8'd8,  9'd168},{  1'b0, 1'b1,   8'd3,  9'd308},
{  1'b0, 1'b0, 8'd173,    9'd0},{  1'b0, 1'b0, 8'd172,    9'd0},{  1'b0, 1'b0, 8'd113,    9'd0},{  1'b0, 1'b0, 8'd104,  9'd345},{  1'b0, 1'b0,  8'd62,  9'd117},{  1'b0, 1'b0,  8'd53,    9'd0},{  1'b0, 1'b0,  8'd43,  9'd319},{  1'b0, 1'b0,  8'd14,  9'd244},{  1'b0, 1'b0,  8'd10,  9'd273},{  1'b0, 1'b1,   8'd6,  9'd123},
{  1'b0, 1'b0, 8'd174,    9'd0},{  1'b0, 1'b0, 8'd173,    9'd0},{  1'b0, 1'b0, 8'd114,    9'd0},{  1'b0, 1'b0,  8'd80,  9'd122},{  1'b0, 1'b0,  8'd70,  9'd249},{  1'b0, 1'b0,  8'd54,    9'd0},{  1'b0, 1'b0,  8'd49,  9'd148},{  1'b0, 1'b0,  8'd17,   9'd66},{  1'b0, 1'b0,  8'd11,  9'd324},{  1'b0, 1'b1,   8'd8,   9'd90},
{  1'b0, 1'b0, 8'd175,    9'd0},{  1'b0, 1'b0, 8'd174,    9'd0},{  1'b0, 1'b0, 8'd118,   9'd94},{  1'b0, 1'b0, 8'd115,    9'd0},{  1'b0, 1'b0, 8'd106,  9'd184},{  1'b0, 1'b0,  8'd55,    9'd0},{  1'b0, 1'b0,  8'd32,  9'd110},{  1'b0, 1'b0,  8'd20,   9'd34},{  1'b0, 1'b0,   8'd8,  9'd177},{  1'b0, 1'b1,   8'd4,  9'd238},
{  1'b0, 1'b0, 8'd176,    9'd0},{  1'b0, 1'b0, 8'd175,    9'd0},{  1'b0, 1'b0, 8'd116,    9'd0},{  1'b0, 1'b0, 8'd109,   9'd58},{  1'b0, 1'b0, 8'd100,   9'd70},{  1'b0, 1'b0,  8'd59,   9'd86},{  1'b0, 1'b0,  8'd56,    9'd0},{  1'b0, 1'b0,  8'd46,  9'd267},{  1'b0, 1'b0,   8'd9,   9'd11},{  1'b0, 1'b1,   8'd2,  9'd242},
{  1'b0, 1'b0, 8'd177,    9'd0},{  1'b0, 1'b0, 8'd176,    9'd0},{  1'b0, 1'b0, 8'd117,    9'd0},{  1'b0, 1'b0,  8'd83,  9'd167},{  1'b0, 1'b0,  8'd63,  9'd223},{  1'b0, 1'b0,  8'd57,    9'd0},{  1'b0, 1'b0,  8'd49,   9'd86},{  1'b0, 1'b0,  8'd43,  9'd183},{  1'b0, 1'b0,  8'd10,   9'd71},{  1'b0, 1'b1,   8'd3,  9'd257},
{  1'b0, 1'b0, 8'd178,    9'd0},{  1'b0, 1'b0, 8'd177,    9'd0},{  1'b0, 1'b0, 8'd118,    9'd0},{  1'b0, 1'b0,  8'd89,   9'd41},{  1'b0, 1'b0,  8'd67,  9'd156},{  1'b0, 1'b0,  8'd58,    9'd0},{  1'b0, 1'b0,  8'd52,   9'd64},{  1'b0, 1'b0,   8'd8,  9'd331},{  1'b0, 1'b0,   8'd5,  9'd162},{  1'b0, 1'b1,   8'd4,   9'd50},
{  1'b0, 1'b0, 8'd179,    9'd0},{  1'b0, 1'b0, 8'd178,    9'd0},{  1'b0, 1'b0, 8'd119,    9'd0},{  1'b0, 1'b0, 8'd110,   9'd23},{  1'b0, 1'b0, 8'd101,  9'd286},{  1'b0, 1'b0,  8'd59,    9'd0},{  1'b0, 1'b0,   8'd8,  9'd245},{  1'b0, 1'b0,   8'd4,   9'd10},{  1'b0, 1'b0,   8'd3,   9'd72},{  1'b0, 1'b1,   8'd1,  9'd296}
};
localparam bit [18 : 0] cLARGE_HS_V_TAB_2BY3_PACKED[cLARGE_HS_TAB_2BY3_PACKED_SIZE] = '{
{8'd179, 1'b0,   10'd0},{8'd179, 1'b1, 10'd590},
{8'd178, 1'b0, 10'd580},{8'd178, 1'b1, 10'd591},
{8'd177, 1'b0, 10'd570},{8'd177, 1'b1, 10'd581},
{8'd176, 1'b0, 10'd560},{8'd176, 1'b1, 10'd571},
{8'd175, 1'b0, 10'd550},{8'd175, 1'b1, 10'd561},
{8'd174, 1'b0, 10'd540},{8'd174, 1'b1, 10'd551},
{8'd173, 1'b0, 10'd530},{8'd173, 1'b1, 10'd541},
{8'd172, 1'b0, 10'd520},{8'd172, 1'b1, 10'd531},
{8'd171, 1'b0, 10'd510},{8'd171, 1'b1, 10'd521},
{8'd170, 1'b0, 10'd500},{8'd170, 1'b1, 10'd511},
{8'd169, 1'b0, 10'd490},{8'd169, 1'b1, 10'd501},
{8'd168, 1'b0, 10'd480},{8'd168, 1'b1, 10'd491},
{8'd167, 1'b0, 10'd470},{8'd167, 1'b1, 10'd481},
{8'd166, 1'b0, 10'd460},{8'd166, 1'b1, 10'd471},
{8'd165, 1'b0, 10'd450},{8'd165, 1'b1, 10'd461},
{8'd164, 1'b0, 10'd440},{8'd164, 1'b1, 10'd451},
{8'd163, 1'b0, 10'd430},{8'd163, 1'b1, 10'd441},
{8'd162, 1'b0, 10'd420},{8'd162, 1'b1, 10'd431},
{8'd161, 1'b0, 10'd410},{8'd161, 1'b1, 10'd421},
{8'd160, 1'b0, 10'd400},{8'd160, 1'b1, 10'd411},
{8'd159, 1'b0, 10'd390},{8'd159, 1'b1, 10'd401},
{8'd158, 1'b0, 10'd380},{8'd158, 1'b1, 10'd391},
{8'd157, 1'b0, 10'd370},{8'd157, 1'b1, 10'd381},
{8'd156, 1'b0, 10'd360},{8'd156, 1'b1, 10'd371},
{8'd155, 1'b0, 10'd350},{8'd155, 1'b1, 10'd361},
{8'd154, 1'b0, 10'd340},{8'd154, 1'b1, 10'd351},
{8'd153, 1'b0, 10'd330},{8'd153, 1'b1, 10'd341},
{8'd152, 1'b0, 10'd320},{8'd152, 1'b1, 10'd331},
{8'd151, 1'b0, 10'd310},{8'd151, 1'b1, 10'd321},
{8'd150, 1'b0, 10'd300},{8'd150, 1'b1, 10'd311},
{8'd149, 1'b0, 10'd290},{8'd149, 1'b1, 10'd301},
{8'd148, 1'b0, 10'd280},{8'd148, 1'b1, 10'd291},
{8'd147, 1'b0, 10'd270},{8'd147, 1'b1, 10'd281},
{8'd146, 1'b0, 10'd260},{8'd146, 1'b1, 10'd271},
{8'd145, 1'b0, 10'd250},{8'd145, 1'b1, 10'd261},
{8'd144, 1'b0, 10'd240},{8'd144, 1'b1, 10'd251},
{8'd143, 1'b0, 10'd230},{8'd143, 1'b1, 10'd241},
{8'd142, 1'b0, 10'd220},{8'd142, 1'b1, 10'd231},
{8'd141, 1'b0, 10'd210},{8'd141, 1'b1, 10'd221},
{8'd140, 1'b0, 10'd200},{8'd140, 1'b1, 10'd211},
{8'd139, 1'b0, 10'd190},{8'd139, 1'b1, 10'd201},
{8'd138, 1'b0, 10'd180},{8'd138, 1'b1, 10'd191},
{8'd137, 1'b0, 10'd170},{8'd137, 1'b1, 10'd181},
{8'd136, 1'b0, 10'd160},{8'd136, 1'b1, 10'd171},
{8'd135, 1'b0, 10'd150},{8'd135, 1'b1, 10'd161},
{8'd134, 1'b0, 10'd140},{8'd134, 1'b1, 10'd151},
{8'd133, 1'b0, 10'd130},{8'd133, 1'b1, 10'd141},
{8'd132, 1'b0, 10'd120},{8'd132, 1'b1, 10'd131},
{8'd131, 1'b0, 10'd110},{8'd131, 1'b1, 10'd121},
{8'd130, 1'b0, 10'd100},{8'd130, 1'b1, 10'd111},
{8'd129, 1'b0,  10'd90},{8'd129, 1'b1, 10'd101},
{8'd128, 1'b0,  10'd80},{8'd128, 1'b1,  10'd91},
{8'd127, 1'b0,  10'd70},{8'd127, 1'b1,  10'd81},
{8'd126, 1'b0,  10'd60},{8'd126, 1'b1,  10'd71},
{8'd125, 1'b0,  10'd50},{8'd125, 1'b1,  10'd61},
{8'd124, 1'b0,  10'd40},{8'd124, 1'b1,  10'd51},
{8'd123, 1'b0,  10'd30},{8'd123, 1'b1,  10'd41},
{8'd122, 1'b0,  10'd20},{8'd122, 1'b1,  10'd31},
{8'd121, 1'b0,  10'd10},{8'd121, 1'b1,  10'd21},
{8'd120, 1'b0,   10'd1},{8'd120, 1'b1,  10'd11},
{8'd119, 1'b0, 10'd492},{8'd119, 1'b0, 10'd502},{8'd119, 1'b1, 10'd592},
{8'd118, 1'b0, 10'd402},{8'd118, 1'b0, 10'd552},{8'd118, 1'b1, 10'd582},
{8'd117, 1'b0,  10'd22},{8'd117, 1'b0, 10'd312},{8'd117, 1'b1, 10'd572},
{8'd116, 1'b0, 10'd482},{8'd116, 1'b0, 10'd512},{8'd116, 1'b1, 10'd562},
{8'd115, 1'b0, 10'd232},{8'd115, 1'b0, 10'd233},{8'd115, 1'b1, 10'd553},
{8'd114, 1'b0,  10'd32},{8'd114, 1'b0, 10'd472},{8'd114, 1'b1, 10'd542},
{8'd113, 1'b0, 10'd282},{8'd113, 1'b0, 10'd332},{8'd113, 1'b1, 10'd532},
{8'd112, 1'b0,  10'd12},{8'd112, 1'b0, 10'd503},{8'd112, 1'b1, 10'd522},
{8'd111, 1'b0,  10'd13},{8'd111, 1'b0, 10'd392},{8'd111, 1'b1, 10'd513},
{8'd110, 1'b0,  10'd82},{8'd110, 1'b0, 10'd504},{8'd110, 1'b1, 10'd593},
{8'd109, 1'b0, 10'd432},{8'd109, 1'b0, 10'd493},{8'd109, 1'b1, 10'd563},
{8'd108, 1'b0, 10'd172},{8'd108, 1'b0, 10'd352},{8'd108, 1'b1, 10'd483},
{8'd107, 1'b0,  10'd83},{8'd107, 1'b0, 10'd152},{8'd107, 1'b1, 10'd473},
{8'd106, 1'b0,  10'd33},{8'd106, 1'b0, 10'd462},{8'd106, 1'b1, 10'd554},
{8'd105, 1'b0, 10'd252},{8'd105, 1'b0, 10'd283},{8'd105, 1'b1, 10'd452},
{8'd104, 1'b0, 10'd333},{8'd104, 1'b0, 10'd442},{8'd104, 1'b1, 10'd533},
{8'd103, 1'b0,  10'd92},{8'd103, 1'b0, 10'd122},{8'd103, 1'b1, 10'd433},
{8'd102, 1'b0, 10'd162},{8'd102, 1'b0, 10'd382},{8'd102, 1'b1, 10'd422},
{8'd101, 1'b0, 10'd412},{8'd101, 1'b0, 10'd523},{8'd101, 1'b1, 10'd594},
{8'd100, 1'b0, 10'd313},{8'd100, 1'b0, 10'd403},{8'd100, 1'b1, 10'd564},
{ 8'd99, 1'b0,  10'd72},{ 8'd99, 1'b0, 10'd372},{ 8'd99, 1'b1, 10'd393},
{ 8'd98, 1'b0, 10'd253},{ 8'd98, 1'b0, 10'd373},{ 8'd98, 1'b1, 10'd383},
{ 8'd97, 1'b0, 10'd112},{ 8'd97, 1'b0, 10'd302},{ 8'd97, 1'b1, 10'd374},
{ 8'd96, 1'b0, 10'd272},{ 8'd96, 1'b0, 10'd362},{ 8'd96, 1'b1, 10'd434},
{ 8'd95, 1'b0, 10'd353},{ 8'd95, 1'b0, 10'd404},{ 8'd95, 1'b1, 10'd524},
{ 8'd94, 1'b0,  10'd93},{ 8'd94, 1'b0, 10'd102},{ 8'd94, 1'b1, 10'd342},
{ 8'd93, 1'b0, 10'd334},{ 8'd93, 1'b0, 10'd394},{ 8'd93, 1'b1, 10'd443},
{ 8'd92, 1'b0, 10'd322},{ 8'd92, 1'b0, 10'd384},{ 8'd92, 1'b1, 10'd484},
{ 8'd91, 1'b0, 10'd292},{ 8'd91, 1'b0, 10'd314},{ 8'd91, 1'b1, 10'd363},
{ 8'd90, 1'b0, 10'd202},{ 8'd90, 1'b0, 10'd303},{ 8'd90, 1'b1, 10'd444},
{ 8'd89, 1'b0, 10'd242},{ 8'd89, 1'b0, 10'd293},{ 8'd89, 1'b1, 10'd583},
{ 8'd88, 1'b0,  10'd73},{ 8'd88, 1'b0, 10'd182},{ 8'd88, 1'b1, 10'd284},
{ 8'd87, 1'b0, 10'd212},{ 8'd87, 1'b0, 10'd273},{ 8'd87, 1'b1, 10'd413},
{ 8'd86, 1'b0, 10'd163},{ 8'd86, 1'b0, 10'd262},{ 8'd86, 1'b1, 10'd304},
{ 8'd85, 1'b0,  10'd23},{ 8'd85, 1'b0, 10'd103},{ 8'd85, 1'b1, 10'd254},
{ 8'd84, 1'b0, 10'd192},{ 8'd84, 1'b0, 10'd243},{ 8'd84, 1'b1, 10'd453},
{ 8'd83, 1'b0,  10'd62},{ 8'd83, 1'b0, 10'd234},{ 8'd83, 1'b1, 10'd573},
{ 8'd82, 1'b0, 10'd113},{ 8'd82, 1'b0, 10'd142},{ 8'd82, 1'b1, 10'd222},
{ 8'd81, 1'b0, 10'd213},{ 8'd81, 1'b0, 10'd214},{ 8'd81, 1'b1, 10'd263},
{ 8'd80, 1'b0, 10'd203},{ 8'd80, 1'b0, 10'd323},{ 8'd80, 1'b1, 10'd543},
{ 8'd79, 1'b0,   10'd2},{ 8'd79, 1'b0,   10'd3},{ 8'd79, 1'b1, 10'd193},
{ 8'd78, 1'b0,  10'd42},{ 8'd78, 1'b0, 10'd173},{ 8'd78, 1'b1, 10'd183},
{ 8'd77, 1'b0, 10'd143},{ 8'd77, 1'b0, 10'd174},{ 8'd77, 1'b1, 10'd264},
{ 8'd76, 1'b0, 10'd132},{ 8'd76, 1'b0, 10'd164},{ 8'd76, 1'b1, 10'd454},
{ 8'd75, 1'b0, 10'd153},{ 8'd75, 1'b0, 10'd423},{ 8'd75, 1'b1, 10'd494},
{ 8'd74, 1'b0, 10'd144},{ 8'd74, 1'b0, 10'd223},{ 8'd74, 1'b1, 10'd514},
{ 8'd73, 1'b0, 10'd133},{ 8'd73, 1'b0, 10'd294},{ 8'd73, 1'b1, 10'd324},
{ 8'd72, 1'b0,  10'd43},{ 8'd72, 1'b0, 10'd123},{ 8'd72, 1'b1, 10'd274},
{ 8'd71, 1'b0, 10'd114},{ 8'd71, 1'b0, 10'd154},{ 8'd71, 1'b1, 10'd364},
{ 8'd70, 1'b0, 10'd104},{ 8'd70, 1'b0, 10'd224},{ 8'd70, 1'b1, 10'd544},
{ 8'd69, 1'b0,  10'd63},{ 8'd69, 1'b0,  10'd94},{ 8'd69, 1'b1, 10'd343},
{ 8'd68, 1'b0,  10'd84},{ 8'd68, 1'b0, 10'd244},{ 8'd68, 1'b1, 10'd354},
{ 8'd67, 1'b0,  10'd74},{ 8'd67, 1'b0, 10'd194},{ 8'd67, 1'b1, 10'd584},
{ 8'd66, 1'b0,  10'd52},{ 8'd66, 1'b0,  10'd64},{ 8'd66, 1'b1, 10'd184},
{ 8'd65, 1'b0,  10'd53},{ 8'd65, 1'b0, 10'd134},{ 8'd65, 1'b1, 10'd344},
{ 8'd64, 1'b0,  10'd44},{ 8'd64, 1'b0, 10'd414},{ 8'd64, 1'b1, 10'd424},
{ 8'd63, 1'b0,  10'd34},{ 8'd63, 1'b0, 10'd124},{ 8'd63, 1'b1, 10'd574},
{ 8'd62, 1'b0,  10'd24},{ 8'd62, 1'b0,  10'd54},{ 8'd62, 1'b1, 10'd534},
{ 8'd61, 1'b0,  10'd14},{ 8'd61, 1'b0, 10'd204},{ 8'd61, 1'b1, 10'd463},
{ 8'd60, 1'b0,   10'd4},{ 8'd60, 1'b0, 10'd464},{ 8'd60, 1'b1, 10'd474},
{ 8'd59, 1'b0, 10'd445},{ 8'd59, 1'b0, 10'd565},{ 8'd59, 1'b1, 10'd595},
{ 8'd58, 1'b0,  10'd45},{ 8'd58, 1'b0, 10'd275},{ 8'd58, 1'b1, 10'd585},
{ 8'd57, 1'b0,  10'd55},{ 8'd57, 1'b0, 10'd345},{ 8'd57, 1'b1, 10'd575},
{ 8'd56, 1'b0, 10'd125},{ 8'd56, 1'b0, 10'd155},{ 8'd56, 1'b1, 10'd566},
{ 8'd55, 1'b0, 10'd225},{ 8'd55, 1'b0, 10'd295},{ 8'd55, 1'b1, 10'd555},
{ 8'd54, 1'b0, 10'd265},{ 8'd54, 1'b0, 10'd266},{ 8'd54, 1'b1, 10'd545},
{ 8'd53, 1'b0, 10'd235},{ 8'd53, 1'b0, 10'd405},{ 8'd53, 1'b1, 10'd535},
{ 8'd52, 1'b0, 10'd346},{ 8'd52, 1'b0, 10'd525},{ 8'd52, 1'b1, 10'd586},
{ 8'd51, 1'b0, 10'd365},{ 8'd51, 1'b0, 10'd515},{ 8'd51, 1'b1, 10'd526},
{ 8'd50, 1'b0, 10'd195},{ 8'd50, 1'b0, 10'd475},{ 8'd50, 1'b1, 10'd505},
{ 8'd49, 1'b0, 10'd495},{ 8'd49, 1'b0, 10'd546},{ 8'd49, 1'b1, 10'd576},
{ 8'd48, 1'b0, 10'd226},{ 8'd48, 1'b0, 10'd425},{ 8'd48, 1'b1, 10'd485},
{ 8'd47, 1'b0,  10'd25},{ 8'd47, 1'b0, 10'd196},{ 8'd47, 1'b1, 10'd476},
{ 8'd46, 1'b0, 10'd415},{ 8'd46, 1'b0, 10'd465},{ 8'd46, 1'b1, 10'd567},
{ 8'd45, 1'b0, 10'd245},{ 8'd45, 1'b0, 10'd455},{ 8'd45, 1'b1, 10'd486},
{ 8'd44, 1'b0, 10'd126},{ 8'd44, 1'b0, 10'd205},{ 8'd44, 1'b1, 10'd446},
{ 8'd43, 1'b0, 10'd435},{ 8'd43, 1'b0, 10'd536},{ 8'd43, 1'b1, 10'd577},
{ 8'd42, 1'b0,  10'd95},{ 8'd42, 1'b0, 10'd105},{ 8'd42, 1'b1, 10'd426},
{ 8'd41, 1'b0, 10'd416},{ 8'd41, 1'b0, 10'd456},{ 8'd41, 1'b1, 10'd466},
{ 8'd40, 1'b0, 10'd135},{ 8'd40, 1'b0, 10'd406},{ 8'd40, 1'b1, 10'd527},
{ 8'd39, 1'b0,   10'd5},{ 8'd39, 1'b0,  10'd26},{ 8'd39, 1'b1, 10'd395},
{ 8'd38, 1'b0, 10'd106},{ 8'd38, 1'b0, 10'd185},{ 8'd38, 1'b1, 10'd385},
{ 8'd37, 1'b0, 10'd255},{ 8'd37, 1'b0, 10'd375},{ 8'd37, 1'b1, 10'd396},
{ 8'd36, 1'b0, 10'd215},{ 8'd36, 1'b0, 10'd366},{ 8'd36, 1'b1, 10'd457},
{ 8'd35, 1'b0,  10'd65},{ 8'd35, 1'b0, 10'd305},{ 8'd35, 1'b1, 10'd355},
{ 8'd34, 1'b0, 10'd165},{ 8'd34, 1'b0, 10'd175},{ 8'd34, 1'b1, 10'd347},
{ 8'd33, 1'b0, 10'd115},{ 8'd33, 1'b0, 10'd335},{ 8'd33, 1'b1, 10'd436},
{ 8'd32, 1'b0, 10'd325},{ 8'd32, 1'b0, 10'd386},{ 8'd32, 1'b1, 10'd556},
{ 8'd31, 1'b0,  10'd85},{ 8'd31, 1'b0, 10'd315},{ 8'd31, 1'b1, 10'd506},
{ 8'd30, 1'b0,  10'd46},{ 8'd30, 1'b0, 10'd276},{ 8'd30, 1'b1, 10'd306},
{ 8'd29, 1'b0, 10'd186},{ 8'd29, 1'b0, 10'd296},{ 8'd29, 1'b1, 10'd397},
{ 8'd28, 1'b0, 10'd216},{ 8'd28, 1'b0, 10'd285},{ 8'd28, 1'b1, 10'd297},
{ 8'd27, 1'b0, 10'd145},{ 8'd27, 1'b0, 10'd277},{ 8'd27, 1'b1, 10'd437},
{ 8'd26, 1'b0, 10'd267},{ 8'd26, 1'b0, 10'd336},{ 8'd26, 1'b1, 10'd356},
{ 8'd25, 1'b0, 10'd156},{ 8'd25, 1'b0, 10'd256},{ 8'd25, 1'b1, 10'd447},
{ 8'd24, 1'b0, 10'd246},{ 8'd24, 1'b0, 10'd417},{ 8'd24, 1'b1, 10'd507},
{ 8'd23, 1'b0, 10'd146},{ 8'd23, 1'b0, 10'd236},{ 8'd23, 1'b1, 10'd357},
{ 8'd22, 1'b0, 10'd227},{ 8'd22, 1'b0, 10'd286},{ 8'd22, 1'b1, 10'd407},
{ 8'd21, 1'b0, 10'd217},{ 8'd21, 1'b0, 10'd387},{ 8'd21, 1'b1, 10'd496},
{ 8'd20, 1'b0, 10'd206},{ 8'd20, 1'b0, 10'd376},{ 8'd20, 1'b1, 10'd557},
{ 8'd19, 1'b0, 10'd166},{ 8'd19, 1'b0, 10'd197},{ 8'd19, 1'b1, 10'd367},
{ 8'd18, 1'b0, 10'd187},{ 8'd18, 1'b0, 10'd307},{ 8'd18, 1'b1, 10'd487},
{ 8'd17, 1'b0,  10'd15},{ 8'd17, 1'b0, 10'd176},{ 8'd17, 1'b1, 10'd547},
{ 8'd16, 1'b0,  10'd35},{ 8'd16, 1'b0, 10'd167},{ 8'd16, 1'b1, 10'd207},
{ 8'd15, 1'b0, 10'd157},{ 8'd15, 1'b0, 10'd427},{ 8'd15, 1'b1, 10'd467},
{ 8'd14, 1'b0,  10'd75},{ 8'd14, 1'b0, 10'd147},{ 8'd14, 1'b1, 10'd537},
{ 8'd13, 1'b0,  10'd86},{ 8'd13, 1'b0, 10'd136},{ 8'd13, 1'b1, 10'd477},
{ 8'd12, 1'b0,   10'd6},{ 8'd12, 1'b0,  10'd16},{ 8'd12, 1'b1, 10'd127},
{ 8'd11, 1'b0,   10'd7},{ 8'd11, 1'b0,  10'd27},{ 8'd11, 1'b0,  10'd87},{ 8'd11, 1'b0, 10'd116},{ 8'd11, 1'b0, 10'd137},{ 8'd11, 1'b0, 10'd237},{ 8'd11, 1'b0, 10'd247},{ 8'd11, 1'b0, 10'd298},{ 8'd11, 1'b0, 10'd316},{ 8'd11, 1'b0, 10'd326},{ 8'd11, 1'b0, 10'd358},{ 8'd11, 1'b0, 10'd398},{ 8'd11, 1'b1, 10'd548},
{ 8'd10, 1'b0,  10'd88},{ 8'd10, 1'b0, 10'd107},{ 8'd10, 1'b0, 10'd158},{ 8'd10, 1'b0, 10'd168},{ 8'd10, 1'b0, 10'd287},{ 8'd10, 1'b0, 10'd288},{ 8'd10, 1'b0, 10'd337},{ 8'd10, 1'b0, 10'd428},{ 8'd10, 1'b0, 10'd458},{ 8'd10, 1'b0, 10'd497},{ 8'd10, 1'b0, 10'd516},{ 8'd10, 1'b0, 10'd538},{ 8'd10, 1'b1, 10'd578},
{  8'd9, 1'b0,  10'd56},{  8'd9, 1'b0,  10'd96},{  8'd9, 1'b0, 10'd128},{  8'd9, 1'b0, 10'd188},{  8'd9, 1'b0, 10'd198},{  8'd9, 1'b0, 10'd257},{  8'd9, 1'b0, 10'd299},{  8'd9, 1'b0, 10'd308},{  8'd9, 1'b0, 10'd338},{  8'd9, 1'b0, 10'd377},{  8'd9, 1'b0, 10'd388},{  8'd9, 1'b0, 10'd438},{  8'd9, 1'b1, 10'd568},
{  8'd8, 1'b0,  10'd28},{  8'd8, 1'b0,  10'd66},{  8'd8, 1'b0,  10'd89},{  8'd8, 1'b0, 10'd117},{  8'd8, 1'b0, 10'd228},{  8'd8, 1'b0, 10'd248},{  8'd8, 1'b0, 10'd468},{  8'd8, 1'b0, 10'd508},{  8'd8, 1'b0, 10'd528},{  8'd8, 1'b0, 10'd549},{  8'd8, 1'b0, 10'd558},{  8'd8, 1'b0, 10'd587},{  8'd8, 1'b1, 10'd596},
{  8'd7, 1'b0,  10'd17},{  8'd7, 1'b0,  10'd57},{  8'd7, 1'b0,  10'd76},{  8'd7, 1'b0,  10'd77},{  8'd7, 1'b0,  10'd97},{  8'd7, 1'b0, 10'd108},{  8'd7, 1'b0, 10'd218},{  8'd7, 1'b0, 10'd219},{  8'd7, 1'b0, 10'd317},{  8'd7, 1'b0, 10'd327},{  8'd7, 1'b0, 10'd348},{  8'd7, 1'b0, 10'd408},{  8'd7, 1'b1, 10'd418},
{  8'd6, 1'b0,  10'd36},{  8'd6, 1'b0,  10'd67},{  8'd6, 1'b0,  10'd68},{  8'd6, 1'b0, 10'd109},{  8'd6, 1'b0, 10'd118},{  8'd6, 1'b0, 10'd177},{  8'd6, 1'b0, 10'd318},{  8'd6, 1'b0, 10'd439},{  8'd6, 1'b0, 10'd459},{  8'd6, 1'b0, 10'd478},{  8'd6, 1'b0, 10'd479},{  8'd6, 1'b0, 10'd517},{  8'd6, 1'b1, 10'd539},
{  8'd5, 1'b0,  10'd58},{  8'd5, 1'b0,  10'd59},{  8'd5, 1'b0,  10'd98},{  8'd5, 1'b0, 10'd178},{  8'd5, 1'b0, 10'd189},{  8'd5, 1'b0, 10'd208},{  8'd5, 1'b0, 10'd309},{  8'd5, 1'b0, 10'd328},{  8'd5, 1'b0, 10'd368},{  8'd5, 1'b0, 10'd429},{  8'd5, 1'b0, 10'd498},{  8'd5, 1'b0, 10'd518},{  8'd5, 1'b1, 10'd588},
{  8'd4, 1'b0,  10'd47},{  8'd4, 1'b0,  10'd99},{  8'd4, 1'b0, 10'd148},{  8'd4, 1'b0, 10'd238},{  8'd4, 1'b0, 10'd268},{  8'd4, 1'b0, 10'd278},{  8'd4, 1'b0, 10'd319},{  8'd4, 1'b0, 10'd389},{  8'd4, 1'b0, 10'd448},{  8'd4, 1'b0, 10'd488},{  8'd4, 1'b0, 10'd559},{  8'd4, 1'b0, 10'd589},{  8'd4, 1'b1, 10'd597},
{  8'd3, 1'b0,  10'd18},{  8'd3, 1'b0,  10'd37},{  8'd3, 1'b0,  10'd38},{  8'd3, 1'b0, 10'd129},{  8'd3, 1'b0, 10'd169},{  8'd3, 1'b0, 10'd229},{  8'd3, 1'b0, 10'd349},{  8'd3, 1'b0, 10'd369},{  8'd3, 1'b0, 10'd378},{  8'd3, 1'b0, 10'd499},{  8'd3, 1'b0, 10'd529},{  8'd3, 1'b0, 10'd579},{  8'd3, 1'b1, 10'd598},
{  8'd2, 1'b0,  10'd29},{  8'd2, 1'b0,  10'd48},{  8'd2, 1'b0, 10'd119},{  8'd2, 1'b0, 10'd149},{  8'd2, 1'b0, 10'd159},{  8'd2, 1'b0, 10'd179},{  8'd2, 1'b0, 10'd249},{  8'd2, 1'b0, 10'd289},{  8'd2, 1'b0, 10'd359},{  8'd2, 1'b0, 10'd379},{  8'd2, 1'b0, 10'd419},{  8'd2, 1'b0, 10'd509},{  8'd2, 1'b1, 10'd569},
{  8'd1, 1'b0,  10'd19},{  8'd1, 1'b0,  10'd39},{  8'd1, 1'b0,  10'd49},{  8'd1, 1'b0,  10'd78},{  8'd1, 1'b0, 10'd138},{  8'd1, 1'b0, 10'd209},{  8'd1, 1'b0, 10'd258},{  8'd1, 1'b0, 10'd279},{  8'd1, 1'b0, 10'd329},{  8'd1, 1'b0, 10'd339},{  8'd1, 1'b0, 10'd409},{  8'd1, 1'b0, 10'd449},{  8'd1, 1'b1, 10'd599},
{  8'd0, 1'b0,   10'd8},{  8'd0, 1'b0,   10'd9},{  8'd0, 1'b0,  10'd69},{  8'd0, 1'b0,  10'd79},{  8'd0, 1'b0, 10'd139},{  8'd0, 1'b0, 10'd199},{  8'd0, 1'b0, 10'd239},{  8'd0, 1'b0, 10'd259},{  8'd0, 1'b0, 10'd269},{  8'd0, 1'b0, 10'd399},{  8'd0, 1'b0, 10'd469},{  8'd0, 1'b0, 10'd489},{  8'd0, 1'b1, 10'd519}
};
localparam int          cLARGE_HS_TAB_3BY4_PACKED_SIZE = 630;
localparam bit [18 : 0] cLARGE_HS_TAB_3BY4_PACKED[cLARGE_HS_TAB_3BY4_PACKED_SIZE] = '{
{  1'b1, 1'b0, 8'd179,    9'd1},{  1'b0, 1'b0, 8'd135,    9'd0},{  1'b0, 1'b0, 8'd126,  9'd282},{  1'b0, 1'b0,  8'd94,  9'd173},{  1'b0, 1'b0,  8'd90,    9'd0},{  1'b0, 1'b0,  8'd69,   9'd59},{  1'b0, 1'b0,  8'd59,  9'd187},{  1'b0, 1'b0,  8'd45,    9'd0},{  1'b0, 1'b0,  8'd31,   9'd97},{  1'b0, 1'b0,  8'd10,  9'd196},{  1'b0, 1'b0,   8'd6,  9'd215},{  1'b0, 1'b0,   8'd3,  9'd155},{  1'b0, 1'b0,   8'd2,  9'd308},{  1'b0, 1'b1,   8'd0,    9'd0},
{  1'b0, 1'b0, 8'd136,    9'd0},{  1'b0, 1'b0, 8'd135,    9'd0},{  1'b0, 1'b0, 8'd129,  9'd180},{  1'b0, 1'b0, 8'd113,  9'd331},{  1'b0, 1'b0,  8'd91,    9'd0},{  1'b0, 1'b0,  8'd82,  9'd209},{  1'b0, 1'b0,  8'd62,  9'd268},{  1'b0, 1'b0,  8'd46,    9'd0},{  1'b0, 1'b0,  8'd40,  9'd181},{  1'b0, 1'b0,  8'd39,  9'd318},{  1'b0, 1'b0,   8'd9,   9'd46},{  1'b0, 1'b0,   8'd7,    9'd9},{  1'b0, 1'b0,   8'd3,   9'd81},{  1'b0, 1'b1,   8'd1,    9'd0},
{  1'b0, 1'b0, 8'd137,    9'd0},{  1'b0, 1'b0, 8'd136,    9'd0},{  1'b0, 1'b0, 8'd114,  9'd332},{  1'b0, 1'b0,  8'd92,    9'd0},{  1'b0, 1'b0,  8'd90,  9'd157},{  1'b0, 1'b0,  8'd85,  9'd327},{  1'b0, 1'b0,  8'd51,  9'd176},{  1'b0, 1'b0,  8'd47,    9'd0},{  1'b0, 1'b0,  8'd40,  9'd347},{  1'b0, 1'b0,  8'd30,   9'd70},{  1'b0, 1'b0,   8'd7,  9'd338},{  1'b0, 1'b0,   8'd2,    9'd0},{  1'b0, 1'b0,   8'd2,  9'd271},{  1'b0, 1'b1,   8'd1,  9'd150},
{  1'b0, 1'b0, 8'd138,    9'd0},{  1'b0, 1'b0, 8'd137,    9'd0},{  1'b0, 1'b0, 8'd134,   9'd64},{  1'b0, 1'b0, 8'd123,  9'd165},{  1'b0, 1'b0,  8'd93,    9'd0},{  1'b0, 1'b0,  8'd50,  9'd155},{  1'b0, 1'b0,  8'd48,    9'd0},{  1'b0, 1'b0,  8'd48,  9'd262},{  1'b0, 1'b0,  8'd17,  9'd291},{  1'b0, 1'b0,   8'd8,   9'd12},{  1'b0, 1'b0,   8'd8,  9'd309},{  1'b0, 1'b0,   8'd7,   9'd88},{  1'b0, 1'b0,   8'd5,  9'd140},{  1'b0, 1'b1,   8'd3,    9'd0},
{  1'b0, 1'b0, 8'd139,    9'd0},{  1'b0, 1'b0, 8'd138,    9'd0},{  1'b0, 1'b0, 8'd107,  9'd189},{  1'b0, 1'b0, 8'd100,   9'd20},{  1'b0, 1'b0,  8'd94,    9'd0},{  1'b0, 1'b0,  8'd49,    9'd0},{  1'b0, 1'b0,  8'd46,  9'd280},{  1'b0, 1'b0,  8'd45,   9'd28},{  1'b0, 1'b0,  8'd36,   9'd41},{  1'b0, 1'b0,  8'd29,  9'd191},{  1'b0, 1'b0,  8'd11,  9'd347},{  1'b0, 1'b0,  8'd10,  9'd157},{  1'b0, 1'b0,   8'd4,    9'd0},{  1'b0, 1'b1,   8'd2,  9'd321},
{  1'b0, 1'b0, 8'd140,    9'd0},{  1'b0, 1'b0, 8'd139,    9'd0},{  1'b0, 1'b0, 8'd131,  9'd336},{  1'b0, 1'b0,  8'd95,    9'd0},{  1'b0, 1'b0,  8'd94,   9'd31},{  1'b0, 1'b0,  8'd77,  9'd269},{  1'b0, 1'b0,  8'd73,  9'd356},{  1'b0, 1'b0,  8'd50,    9'd0},{  1'b0, 1'b0,  8'd32,  9'd305},{  1'b0, 1'b0,  8'd30,   9'd77},{  1'b0, 1'b0,   8'd9,  9'd161},{  1'b0, 1'b0,   8'd5,    9'd0},{  1'b0, 1'b0,   8'd5,  9'd278},{  1'b0, 1'b1,   8'd5,   9'd31},
{  1'b0, 1'b0, 8'd141,    9'd0},{  1'b0, 1'b0, 8'd140,    9'd0},{  1'b0, 1'b0, 8'd106,   9'd61},{  1'b0, 1'b0,  8'd98,  9'd107},{  1'b0, 1'b0,  8'd96,    9'd0},{  1'b0, 1'b0,  8'd89,  9'd138},{  1'b0, 1'b0,  8'd51,    9'd0},{  1'b0, 1'b0,  8'd48,   9'd70},{  1'b0, 1'b0,  8'd16,  9'd298},{  1'b0, 1'b0,  8'd12,  9'd194},{  1'b0, 1'b0,   8'd9,   9'd12},{  1'b0, 1'b0,   8'd8,  9'd204},{  1'b0, 1'b0,   8'd6,    9'd0},{  1'b0, 1'b1,   8'd5,  9'd315},
{  1'b0, 1'b0, 8'd142,    9'd0},{  1'b0, 1'b0, 8'd141,    9'd0},{  1'b0, 1'b0, 8'd123,  9'd299},{  1'b0, 1'b0, 8'd108,  9'd198},{  1'b0, 1'b0,  8'd97,    9'd0},{  1'b0, 1'b0,  8'd66,   9'd87},{  1'b0, 1'b0,  8'd52,    9'd0},{  1'b0, 1'b0,  8'd47,   9'd60},{  1'b0, 1'b0,  8'd33,  9'd315},{  1'b0, 1'b0,  8'd19,  9'd160},{  1'b0, 1'b0,  8'd14,  9'd181},{  1'b0, 1'b0,  8'd13,  9'd150},{  1'b0, 1'b0,   8'd9,  9'd281},{  1'b0, 1'b1,   8'd7,    9'd0},
{  1'b0, 1'b0, 8'd143,    9'd0},{  1'b0, 1'b0, 8'd142,    9'd0},{  1'b0, 1'b0, 8'd116,  9'd146},{  1'b0, 1'b0,  8'd98,    9'd0},{  1'b0, 1'b0,  8'd96,  9'd171},{  1'b0, 1'b0,  8'd89,  9'd171},{  1'b0, 1'b0,  8'd55,   9'd39},{  1'b0, 1'b0,  8'd53,    9'd0},{  1'b0, 1'b0,  8'd21,   9'd98},{  1'b0, 1'b0,  8'd12,  9'd328},{  1'b0, 1'b0,  8'd10,  9'd224},{  1'b0, 1'b0,   8'd8,    9'd0},{  1'b0, 1'b0,   8'd8,   9'd79},{  1'b0, 1'b1,   8'd4,   9'd36},
{  1'b0, 1'b0, 8'd144,    9'd0},{  1'b0, 1'b0, 8'd143,    9'd0},{  1'b0, 1'b0, 8'd111,   9'd89},{  1'b0, 1'b0, 8'd108,  9'd271},{  1'b0, 1'b0,  8'd99,    9'd0},{  1'b0, 1'b0,  8'd87,   9'd26},{  1'b0, 1'b0,  8'd57,   9'd12},{  1'b0, 1'b0,  8'd54,    9'd0},{  1'b0, 1'b0,  8'd29,  9'd285},{  1'b0, 1'b0,   8'd9,    9'd0},{  1'b0, 1'b0,   8'd6,   9'd90},{  1'b0, 1'b0,   8'd4,  9'd240},{  1'b0, 1'b0,   8'd2,  9'd142},{  1'b0, 1'b1,   8'd1,  9'd307},
{  1'b0, 1'b0, 8'd145,    9'd0},{  1'b0, 1'b0, 8'd144,    9'd0},{  1'b0, 1'b0, 8'd100,    9'd0},{  1'b0, 1'b0, 8'd100,   9'd40},{  1'b0, 1'b0,  8'd99,  9'd265},{  1'b0, 1'b0,  8'd78,  9'd344},{  1'b0, 1'b0,  8'd63,  9'd179},{  1'b0, 1'b0,  8'd55,    9'd0},{  1'b0, 1'b0,  8'd13,   9'd11},{  1'b0, 1'b0,  8'd12,   9'd81},{  1'b0, 1'b0,  8'd10,    9'd0},{  1'b0, 1'b0,   8'd9,  9'd147},{  1'b0, 1'b0,   8'd4,  9'd108},{  1'b0, 1'b1,   8'd1,  9'd340},
{  1'b0, 1'b0, 8'd146,    9'd0},{  1'b0, 1'b0, 8'd145,    9'd0},{  1'b0, 1'b0, 8'd122,  9'd272},{  1'b0, 1'b0, 8'd101,    9'd0},{  1'b0, 1'b0,  8'd97,   9'd57},{  1'b0, 1'b0,  8'd57,  9'd276},{  1'b0, 1'b0,  8'd56,    9'd0},{  1'b0, 1'b0,  8'd56,   9'd38},{  1'b0, 1'b0,  8'd23,  9'd168},{  1'b0, 1'b0,  8'd15,  9'd266},{  1'b0, 1'b0,  8'd11,    9'd0},{  1'b0, 1'b0,   8'd8,  9'd128},{  1'b0, 1'b0,   8'd5,  9'd120},{  1'b0, 1'b1,   8'd0,   9'd18},
{  1'b0, 1'b0, 8'd147,    9'd0},{  1'b0, 1'b0, 8'd146,    9'd0},{  1'b0, 1'b0, 8'd104,  9'd174},{  1'b0, 1'b0, 8'd102,    9'd0},{  1'b0, 1'b0,  8'd90,   9'd77},{  1'b0, 1'b0,  8'd76,  9'd213},{  1'b0, 1'b0,  8'd57,    9'd0},{  1'b0, 1'b0,  8'd52,  9'd335},{  1'b0, 1'b0,  8'd31,  9'd309},{  1'b0, 1'b0,  8'd13,   9'd58},{  1'b0, 1'b0,  8'd12,    9'd0},{  1'b0, 1'b0,  8'd12,  9'd109},{  1'b0, 1'b0,   8'd2,  9'd177},{  1'b0, 1'b1,   8'd0,   9'd72},
{  1'b0, 1'b0, 8'd148,    9'd0},{  1'b0, 1'b0, 8'd147,    9'd0},{  1'b0, 1'b0, 8'd110,  9'd280},{  1'b0, 1'b0, 8'd107,  9'd103},{  1'b0, 1'b0, 8'd103,    9'd0},{  1'b0, 1'b0,  8'd68,   9'd39},{  1'b0, 1'b0,  8'd58,    9'd0},{  1'b0, 1'b0,  8'd53,  9'd112},{  1'b0, 1'b0,  8'd41,  9'd249},{  1'b0, 1'b0,  8'd13,    9'd0},{  1'b0, 1'b0,  8'd13,  9'd198},{  1'b0, 1'b0,  8'd11,   9'd42},{  1'b0, 1'b0,  8'd10,  9'd205},{  1'b0, 1'b1,   8'd4,  9'd206},
{  1'b0, 1'b0, 8'd149,    9'd0},{  1'b0, 1'b0, 8'd148,    9'd0},{  1'b0, 1'b0, 8'd116,  9'd190},{  1'b0, 1'b0, 8'd105,  9'd135},{  1'b0, 1'b0, 8'd104,    9'd0},{  1'b0, 1'b0,  8'd62,   9'd31},{  1'b0, 1'b0,  8'd59,    9'd0},{  1'b0, 1'b0,  8'd51,  9'd357},{  1'b0, 1'b0,  8'd22,   9'd59},{  1'b0, 1'b0,  8'd14,    9'd0},{  1'b0, 1'b0,  8'd13,  9'd294},{  1'b0, 1'b0,  8'd12,  9'd354},{  1'b0, 1'b0,   8'd4,  9'd215},{  1'b0, 1'b1,   8'd3,  9'd262},
{  1'b0, 1'b0, 8'd150,    9'd0},{  1'b0, 1'b0, 8'd149,    9'd0},{  1'b0, 1'b0, 8'd125,   9'd56},{  1'b0, 1'b0, 8'd105,    9'd0},{  1'b0, 1'b0, 8'd102,   9'd79},{  1'b0, 1'b0,  8'd86,  9'd341},{  1'b0, 1'b0,  8'd68,  9'd130},{  1'b0, 1'b0,  8'd60,    9'd0},{  1'b0, 1'b0,  8'd26,  9'd136},{  1'b0, 1'b0,  8'd18,  9'd321},{  1'b0, 1'b0,  8'd15,    9'd0},{  1'b0, 1'b0,  8'd10,  9'd146},{  1'b0, 1'b0,   8'd7,  9'd267},{  1'b0, 1'b1,   8'd4,   9'd27},
{  1'b0, 1'b0, 8'd151,    9'd0},{  1'b0, 1'b0, 8'd150,    9'd0},{  1'b0, 1'b0, 8'd114,  9'd158},{  1'b0, 1'b0, 8'd106,    9'd0},{  1'b0, 1'b0,  8'd91,   9'd87},{  1'b0, 1'b0,  8'd85,  9'd188},{  1'b0, 1'b0,  8'd84,  9'd189},{  1'b0, 1'b0,  8'd61,    9'd0},{  1'b0, 1'b0,  8'd35,  9'd117},{  1'b0, 1'b0,  8'd16,    9'd0},{  1'b0, 1'b0,   8'd9,  9'd217},{  1'b0, 1'b0,   8'd6,  9'd196},{  1'b0, 1'b0,   8'd6,  9'd103},{  1'b0, 1'b1,   8'd3,  9'd162},
{  1'b0, 1'b0, 8'd152,    9'd0},{  1'b0, 1'b0, 8'd151,    9'd0},{  1'b0, 1'b0, 8'd129,  9'd226},{  1'b0, 1'b0, 8'd107,    9'd0},{  1'b0, 1'b0, 8'd102,  9'd251},{  1'b0, 1'b0,  8'd88,   9'd52},{  1'b0, 1'b0,  8'd69,  9'd332},{  1'b0, 1'b0,  8'd62,    9'd0},{  1'b0, 1'b0,  8'd39,  9'd170},{  1'b0, 1'b0,  8'd28,  9'd192},{  1'b0, 1'b0,  8'd17,    9'd0},{  1'b0, 1'b0,   8'd3,  9'd295},{  1'b0, 1'b0,   8'd3,  9'd318},{  1'b0, 1'b1,   8'd2,  9'd336},
{  1'b0, 1'b0, 8'd153,    9'd0},{  1'b0, 1'b0, 8'd152,    9'd0},{  1'b0, 1'b0, 8'd121,  9'd255},{  1'b0, 1'b0, 8'd119,  9'd308},{  1'b0, 1'b0, 8'd108,    9'd0},{  1'b0, 1'b0,  8'd63,    9'd0},{  1'b0, 1'b0,  8'd60,  9'd217},{  1'b0, 1'b0,  8'd50,  9'd312},{  1'b0, 1'b0,  8'd18,    9'd0},{  1'b0, 1'b0,  8'd14,  9'd321},{  1'b0, 1'b0,  8'd11,  9'd240},{  1'b0, 1'b0,   8'd7,  9'd203},{  1'b0, 1'b0,   8'd6,  9'd230},{  1'b0, 1'b1,   8'd6,  9'd228},
{  1'b0, 1'b0, 8'd154,    9'd0},{  1'b0, 1'b0, 8'd153,    9'd0},{  1'b0, 1'b0, 8'd127,  9'd207},{  1'b0, 1'b0, 8'd109,    9'd0},{  1'b0, 1'b0,  8'd96,   9'd55},{  1'b0, 1'b0,  8'd87,  9'd176},{  1'b0, 1'b0,  8'd77,  9'd342},{  1'b0, 1'b0,  8'd64,    9'd0},{  1'b0, 1'b0,  8'd35,  9'd334},{  1'b0, 1'b0,  8'd19,    9'd0},{  1'b0, 1'b0,  8'd13,  9'd346},{  1'b0, 1'b0,  8'd12,   9'd47},{  1'b0, 1'b0,   8'd4,  9'd324},{  1'b0, 1'b1,   8'd1,  9'd252},
{  1'b0, 1'b0, 8'd155,    9'd0},{  1'b0, 1'b0, 8'd154,    9'd0},{  1'b0, 1'b0, 8'd132,  9'd321},{  1'b0, 1'b0, 8'd113,   9'd38},{  1'b0, 1'b0, 8'd110,    9'd0},{  1'b0, 1'b0,  8'd74,  9'd103},{  1'b0, 1'b0,  8'd65,    9'd0},{  1'b0, 1'b0,  8'd46,  9'd221},{  1'b0, 1'b0,  8'd38,  9'd135},{  1'b0, 1'b0,  8'd27,  9'd166},{  1'b0, 1'b0,  8'd20,    9'd0},{  1'b0, 1'b0,  8'd10,  9'd246},{  1'b0, 1'b0,   8'd8,   9'd19},{  1'b0, 1'b1,   8'd5,  9'd309},
{  1'b0, 1'b0, 8'd156,    9'd0},{  1'b0, 1'b0, 8'd155,    9'd0},{  1'b0, 1'b0, 8'd111,    9'd0},{  1'b0, 1'b0, 8'd110,   9'd98},{  1'b0, 1'b0, 8'd103,  9'd331},{  1'b0, 1'b0,  8'd82,  9'd106},{  1'b0, 1'b0,  8'd66,    9'd0},{  1'b0, 1'b0,  8'd56,  9'd180},{  1'b0, 1'b0,  8'd21,    9'd0},{  1'b0, 1'b0,  8'd16,  9'd153},{  1'b0, 1'b0,  8'd11,  9'd245},{  1'b0, 1'b0,   8'd4,  9'd169},{  1'b0, 1'b0,   8'd2,  9'd140},{  1'b0, 1'b1,   8'd1,   9'd44},
{  1'b0, 1'b0, 8'd157,    9'd0},{  1'b0, 1'b0, 8'd156,    9'd0},{  1'b0, 1'b0, 8'd120,  9'd263},{  1'b0, 1'b0, 8'd112,    9'd0},{  1'b0, 1'b0,  8'd98,  9'd348},{  1'b0, 1'b0,  8'd84,   9'd62},{  1'b0, 1'b0,  8'd81,  9'd183},{  1'b0, 1'b0,  8'd67,    9'd0},{  1'b0, 1'b0,  8'd22,    9'd0},{  1'b0, 1'b0,   8'd9,  9'd162},{  1'b0, 1'b0,   8'd8,  9'd133},{  1'b0, 1'b0,   8'd4,  9'd253},{  1'b0, 1'b0,   8'd2,  9'd302},{  1'b0, 1'b1,   8'd0,   9'd60},
{  1'b0, 1'b0, 8'd158,    9'd0},{  1'b0, 1'b0, 8'd157,    9'd0},{  1'b0, 1'b0, 8'd113,    9'd0},{  1'b0, 1'b0, 8'd109,  9'd276},{  1'b0, 1'b0, 8'd106,   9'd87},{  1'b0, 1'b0,  8'd68,    9'd0},{  1'b0, 1'b0,  8'd64,  9'd187},{  1'b0, 1'b0,  8'd55,  9'd343},{  1'b0, 1'b0,  8'd36,   9'd24},{  1'b0, 1'b0,  8'd23,    9'd0},{  1'b0, 1'b0,  8'd23,  9'd200},{  1'b0, 1'b0,   8'd6,  9'd174},{  1'b0, 1'b0,   8'd5,  9'd163},{  1'b0, 1'b1,   8'd0,  9'd116},
{  1'b0, 1'b0, 8'd159,    9'd0},{  1'b0, 1'b0, 8'd158,    9'd0},{  1'b0, 1'b0, 8'd133,  9'd247},{  1'b0, 1'b0, 8'd124,  9'd291},{  1'b0, 1'b0, 8'd114,    9'd0},{  1'b0, 1'b0,  8'd80,  9'd345},{  1'b0, 1'b0,  8'd78,  9'd194},{  1'b0, 1'b0,  8'd69,    9'd0},{  1'b0, 1'b0,  8'd38,  9'd214},{  1'b0, 1'b0,  8'd27,  9'd323},{  1'b0, 1'b0,  8'd24,    9'd0},{  1'b0, 1'b0,  8'd11,  9'd328},{  1'b0, 1'b0,   8'd9,   9'd75},{  1'b0, 1'b1,   8'd0,  9'd297},
{  1'b0, 1'b0, 8'd160,    9'd0},{  1'b0, 1'b0, 8'd159,    9'd0},{  1'b0, 1'b0, 8'd118,  9'd284},{  1'b0, 1'b0, 8'd115,    9'd0},{  1'b0, 1'b0,  8'd92,  9'd170},{  1'b0, 1'b0,  8'd81,   9'd66},{  1'b0, 1'b0,  8'd79,  9'd340},{  1'b0, 1'b0,  8'd70,    9'd0},{  1'b0, 1'b0,  8'd42,  9'd303},{  1'b0, 1'b0,  8'd25,    9'd0},{  1'b0, 1'b0,  8'd22,  9'd310},{  1'b0, 1'b0,  8'd11,  9'd256},{  1'b0, 1'b0,   8'd9,  9'd106},{  1'b0, 1'b1,   8'd8,  9'd138},
{  1'b0, 1'b0, 8'd161,    9'd0},{  1'b0, 1'b0, 8'd160,    9'd0},{  1'b0, 1'b0, 8'd128,  9'd341},{  1'b0, 1'b0, 8'd120,  9'd248},{  1'b0, 1'b0, 8'd116,    9'd0},{  1'b0, 1'b0,  8'd71,    9'd0},{  1'b0, 1'b0,  8'd67,   9'd85},{  1'b0, 1'b0,  8'd58,  9'd157},{  1'b0, 1'b0,  8'd26,    9'd0},{  1'b0, 1'b0,  8'd25,  9'd161},{  1'b0, 1'b0,  8'd14,   9'd67},{  1'b0, 1'b0,  8'd14,  9'd145},{  1'b0, 1'b0,   8'd7,  9'd271},{  1'b0, 1'b1,   8'd0,  9'd175},
{  1'b0, 1'b0, 8'd162,    9'd0},{  1'b0, 1'b0, 8'd161,    9'd0},{  1'b0, 1'b0, 8'd118,    9'd6},{  1'b0, 1'b0, 8'd117,    9'd0},{  1'b0, 1'b0,  8'd97,  9'd175},{  1'b0, 1'b0,  8'd73,  9'd169},{  1'b0, 1'b0,  8'd72,    9'd0},{  1'b0, 1'b0,  8'd47,  9'd182},{  1'b0, 1'b0,  8'd34,  9'd292},{  1'b0, 1'b0,  8'd27,    9'd0},{  1'b0, 1'b0,  8'd20,   9'd73},{  1'b0, 1'b0,   8'd9,  9'd109},{  1'b0, 1'b0,   8'd8,  9'd315},{  1'b0, 1'b1,   8'd6,  9'd177},
{  1'b0, 1'b0, 8'd163,    9'd0},{  1'b0, 1'b0, 8'd162,    9'd0},{  1'b0, 1'b0, 8'd128,  9'd311},{  1'b0, 1'b0, 8'd118,    9'd0},{  1'b0, 1'b0, 8'd112,  9'd188},{  1'b0, 1'b0,  8'd75,  9'd291},{  1'b0, 1'b0,  8'd73,    9'd0},{  1'b0, 1'b0,  8'd71,   9'd95},{  1'b0, 1'b0,  8'd43,  9'd190},{  1'b0, 1'b0,  8'd28,    9'd0},{  1'b0, 1'b0,  8'd25,  9'd158},{  1'b0, 1'b0,  8'd14,  9'd349},{  1'b0, 1'b0,  8'd14,  9'd194},{  1'b0, 1'b1,  8'd10,  9'd159},
{  1'b0, 1'b0, 8'd164,    9'd0},{  1'b0, 1'b0, 8'd163,    9'd0},{  1'b0, 1'b0, 8'd119,    9'd0},{  1'b0, 1'b0, 8'd104,  9'd170},{  1'b0, 1'b0,  8'd92,  9'd286},{  1'b0, 1'b0,  8'd80,   9'd64},{  1'b0, 1'b0,  8'd74,    9'd0},{  1'b0, 1'b0,  8'd49,   9'd33},{  1'b0, 1'b0,  8'd29,    9'd0},{  1'b0, 1'b0,  8'd18,   9'd44},{  1'b0, 1'b0,  8'd12,   9'd32},{  1'b0, 1'b0,  8'd11,    9'd2},{  1'b0, 1'b0,   8'd5,  9'd126},{  1'b0, 1'b1,   8'd0,   9'd55},
{  1'b0, 1'b0, 8'd165,    9'd0},{  1'b0, 1'b0, 8'd164,    9'd0},{  1'b0, 1'b0, 8'd126,  9'd143},{  1'b0, 1'b0, 8'd120,    9'd0},{  1'b0, 1'b0,  8'd91,  9'd307},{  1'b0, 1'b0,  8'd75,    9'd0},{  1'b0, 1'b0,  8'd70,  9'd123},{  1'b0, 1'b0,  8'd65,  9'd313},{  1'b0, 1'b0,  8'd30,    9'd0},{  1'b0, 1'b0,  8'd20,   9'd87},{  1'b0, 1'b0,  8'd10,  9'd165},{  1'b0, 1'b0,   8'd6,   9'd75},{  1'b0, 1'b0,   8'd6,  9'd132},{  1'b0, 1'b1,   8'd3,   9'd34},
{  1'b0, 1'b0, 8'd166,    9'd0},{  1'b0, 1'b0, 8'd165,    9'd0},{  1'b0, 1'b0, 8'd134,  9'd322},{  1'b0, 1'b0, 8'd121,    9'd0},{  1'b0, 1'b0,  8'd99,  9'd231},{  1'b0, 1'b0,  8'd76,    9'd0},{  1'b0, 1'b0,  8'd71,  9'd280},{  1'b0, 1'b0,  8'd59,   9'd31},{  1'b0, 1'b0,  8'd44,   9'd59},{  1'b0, 1'b0,  8'd31,    9'd0},{  1'b0, 1'b0,  8'd13,   9'd93},{  1'b0, 1'b0,   8'd7,   9'd98},{  1'b0, 1'b0,   8'd4,  9'd338},{  1'b0, 1'b1,   8'd0,  9'd324},
{  1'b0, 1'b0, 8'd167,    9'd0},{  1'b0, 1'b0, 8'd166,    9'd0},{  1'b0, 1'b0, 8'd127,  9'd152},{  1'b0, 1'b0, 8'd122,    9'd0},{  1'b0, 1'b0, 8'd119,  9'd148},{  1'b0, 1'b0,  8'd77,    9'd0},{  1'b0, 1'b0,  8'd70,  9'd140},{  1'b0, 1'b0,  8'd45,   9'd22},{  1'b0, 1'b0,  8'd32,    9'd0},{  1'b0, 1'b0,  8'd17,  9'd296},{  1'b0, 1'b0,   8'd8,   9'd77},{  1'b0, 1'b0,   8'd3,   9'd84},{  1'b0, 1'b0,   8'd2,  9'd174},{  1'b0, 1'b1,   8'd1,  9'd253},
{  1'b0, 1'b0, 8'd168,    9'd0},{  1'b0, 1'b0, 8'd167,    9'd0},{  1'b0, 1'b0, 8'd130,  9'd107},{  1'b0, 1'b0, 8'd123,    9'd0},{  1'b0, 1'b0,  8'd95,  9'd204},{  1'b0, 1'b0,  8'd78,    9'd0},{  1'b0, 1'b0,  8'd65,   9'd28},{  1'b0, 1'b0,  8'd52,  9'd269},{  1'b0, 1'b0,  8'd42,  9'd138},{  1'b0, 1'b0,  8'd37,   9'd45},{  1'b0, 1'b0,  8'd33,    9'd0},{  1'b0, 1'b0,  8'd14,  9'd248},{  1'b0, 1'b0,  8'd14,  9'd335},{  1'b0, 1'b1,  8'd10,  9'd225},
{  1'b0, 1'b0, 8'd169,    9'd0},{  1'b0, 1'b0, 8'd168,    9'd0},{  1'b0, 1'b0, 8'd124,    9'd0},{  1'b0, 1'b0, 8'd109,  9'd127},{  1'b0, 1'b0, 8'd105,  9'd290},{  1'b0, 1'b0,  8'd79,    9'd0},{  1'b0, 1'b0,  8'd61,  9'd251},{  1'b0, 1'b0,  8'd58,   9'd91},{  1'b0, 1'b0,  8'd37,   9'd23},{  1'b0, 1'b0,  8'd34,    9'd0},{  1'b0, 1'b0,  8'd34,   9'd54},{  1'b0, 1'b0,  8'd12,  9'd352},{  1'b0, 1'b0,   8'd7,  9'd165},{  1'b0, 1'b1,   8'd2,  9'd298},
{  1'b0, 1'b0, 8'd170,    9'd0},{  1'b0, 1'b0, 8'd169,    9'd0},{  1'b0, 1'b0, 8'd125,    9'd0},{  1'b0, 1'b0, 8'd122,  9'd358},{  1'b0, 1'b0, 8'd112,  9'd307},{  1'b0, 1'b0,  8'd86,  9'd173},{  1'b0, 1'b0,  8'd80,    9'd0},{  1'b0, 1'b0,  8'd53,  9'd143},{  1'b0, 1'b0,  8'd35,    9'd0},{  1'b0, 1'b0,  8'd26,  9'd303},{  1'b0, 1'b0,  8'd14,  9'd285},{  1'b0, 1'b0,  8'd11,    9'd4},{  1'b0, 1'b0,   8'd5,   9'd35},{  1'b0, 1'b1,   8'd3,  9'd128},
{  1'b0, 1'b0, 8'd171,    9'd0},{  1'b0, 1'b0, 8'd170,    9'd0},{  1'b0, 1'b0, 8'd126,    9'd0},{  1'b0, 1'b0, 8'd124,  9'd322},{  1'b0, 1'b0, 8'd117,    9'd8},{  1'b0, 1'b0,  8'd81,    9'd0},{  1'b0, 1'b0,  8'd79,  9'd164},{  1'b0, 1'b0,  8'd66,  9'd307},{  1'b0, 1'b0,  8'd36,    9'd0},{  1'b0, 1'b0,  8'd28,   9'd54},{  1'b0, 1'b0,  8'd13,  9'd184},{  1'b0, 1'b0,   8'd6,  9'd340},{  1'b0, 1'b0,   8'd5,  9'd352},{  1'b0, 1'b1,   8'd3,  9'd174},
{  1'b0, 1'b0, 8'd172,    9'd0},{  1'b0, 1'b0, 8'd171,    9'd0},{  1'b0, 1'b0, 8'd133,  9'd114},{  1'b0, 1'b0, 8'd127,    9'd0},{  1'b0, 1'b0, 8'd101,  9'd251},{  1'b0, 1'b0,  8'd82,    9'd0},{  1'b0, 1'b0,  8'd76,  9'd310},{  1'b0, 1'b0,  8'd54,  9'd331},{  1'b0, 1'b0,  8'd37,    9'd0},{  1'b0, 1'b0,  8'd14,  9'd107},{  1'b0, 1'b0,  8'd13,  9'd176},{  1'b0, 1'b0,  8'd12,   9'd59},{  1'b0, 1'b0,   8'd9,   9'd71},{  1'b0, 1'b1,   8'd1,  9'd283},
{  1'b0, 1'b0, 8'd173,    9'd0},{  1'b0, 1'b0, 8'd172,    9'd0},{  1'b0, 1'b0, 8'd130,  9'd265},{  1'b0, 1'b0, 8'd128,    9'd0},{  1'b0, 1'b0, 8'd125,  9'd249},{  1'b0, 1'b0,  8'd88,  9'd192},{  1'b0, 1'b0,  8'd83,    9'd0},{  1'b0, 1'b0,  8'd64,   9'd64},{  1'b0, 1'b0,  8'd38,    9'd0},{  1'b0, 1'b0,  8'd33,  9'd243},{  1'b0, 1'b0,  8'd21,  9'd138},{  1'b0, 1'b0,  8'd14,  9'd303},{  1'b0, 1'b0,  8'd10,   9'd10},{  1'b0, 1'b1,   8'd7,  9'd281},
{  1'b0, 1'b0, 8'd174,    9'd0},{  1'b0, 1'b0, 8'd173,    9'd0},{  1'b0, 1'b0, 8'd129,    9'd0},{  1'b0, 1'b0, 8'd111,   9'd29},{  1'b0, 1'b0, 8'd101,  9'd205},{  1'b0, 1'b0,  8'd84,    9'd0},{  1'b0, 1'b0,  8'd83,  9'd107},{  1'b0, 1'b0,  8'd49,    9'd7},{  1'b0, 1'b0,  8'd39,    9'd0},{  1'b0, 1'b0,  8'd32,  9'd133},{  1'b0, 1'b0,  8'd19,   9'd95},{  1'b0, 1'b0,  8'd10,  9'd291},{  1'b0, 1'b0,   8'd7,   9'd46},{  1'b0, 1'b1,   8'd0,  9'd163},
{  1'b0, 1'b0, 8'd175,    9'd0},{  1'b0, 1'b0, 8'd174,    9'd0},{  1'b0, 1'b0, 8'd130,    9'd0},{  1'b0, 1'b0, 8'd121,  9'd319},{  1'b0, 1'b0, 8'd103,   9'd58},{  1'b0, 1'b0,  8'd85,    9'd0},{  1'b0, 1'b0,  8'd67,   9'd88},{  1'b0, 1'b0,  8'd61,  9'd139},{  1'b0, 1'b0,  8'd40,    9'd0},{  1'b0, 1'b0,  8'd13,   9'd84},{  1'b0, 1'b0,  8'd12,  9'd158},{  1'b0, 1'b0,  8'd11,  9'd235},{  1'b0, 1'b0,   8'd0,  9'd141},{  1'b0, 1'b1,   8'd0,  9'd248},
{  1'b0, 1'b0, 8'd176,    9'd0},{  1'b0, 1'b0, 8'd175,    9'd0},{  1'b0, 1'b0, 8'd132,  9'd178},{  1'b0, 1'b0, 8'd131,    9'd0},{  1'b0, 1'b0,  8'd95,  9'd130},{  1'b0, 1'b0,  8'd86,    9'd0},{  1'b0, 1'b0,  8'd83,  9'd246},{  1'b0, 1'b0,  8'd72,  9'd271},{  1'b0, 1'b0,  8'd44,  9'd260},{  1'b0, 1'b0,  8'd41,    9'd0},{  1'b0, 1'b0,  8'd13,   9'd17},{  1'b0, 1'b0,  8'd11,  9'd176},{  1'b0, 1'b0,   8'd8,  9'd186},{  1'b0, 1'b1,   8'd5,  9'd209},
{  1'b0, 1'b0, 8'd177,    9'd0},{  1'b0, 1'b0, 8'd176,    9'd0},{  1'b0, 1'b0, 8'd132,    9'd0},{  1'b0, 1'b0, 8'd117,  9'd109},{  1'b0, 1'b0,  8'd93,  9'd181},{  1'b0, 1'b0,  8'd87,    9'd0},{  1'b0, 1'b0,  8'd63,  9'd201},{  1'b0, 1'b0,  8'd54,  9'd281},{  1'b0, 1'b0,  8'd42,    9'd0},{  1'b0, 1'b0,  8'd24,  9'd314},{  1'b0, 1'b0,  8'd24,   9'd65},{  1'b0, 1'b0,   8'd3,  9'd194},{  1'b0, 1'b0,   8'd1,    9'd7},{  1'b0, 1'b1,   8'd1,   9'd18},
{  1'b0, 1'b0, 8'd178,    9'd0},{  1'b0, 1'b0, 8'd177,    9'd0},{  1'b0, 1'b0, 8'd133,    9'd0},{  1'b0, 1'b0, 8'd115,  9'd332},{  1'b0, 1'b0, 8'd115,  9'd196},{  1'b0, 1'b0,  8'd88,    9'd0},{  1'b0, 1'b0,  8'd74,  9'd313},{  1'b0, 1'b0,  8'd72,  9'd258},{  1'b0, 1'b0,  8'd43,    9'd0},{  1'b0, 1'b0,  8'd41,  9'd101},{  1'b0, 1'b0,  8'd11,  9'd167},{  1'b0, 1'b0,   8'd4,   9'd46},{  1'b0, 1'b0,   8'd2,   9'd37},{  1'b0, 1'b1,   8'd1,   9'd59},
{  1'b0, 1'b0, 8'd179,    9'd0},{  1'b0, 1'b0, 8'd178,    9'd0},{  1'b0, 1'b0, 8'd134,    9'd0},{  1'b0, 1'b0, 8'd131,  9'd135},{  1'b0, 1'b0,  8'd93,   9'd38},{  1'b0, 1'b0,  8'd89,    9'd0},{  1'b0, 1'b0,  8'd75,  9'd212},{  1'b0, 1'b0,  8'd60,  9'd168},{  1'b0, 1'b0,  8'd44,    9'd0},{  1'b0, 1'b0,  8'd43,  9'd174},{  1'b0, 1'b0,  8'd15,   9'd69},{  1'b0, 1'b0,  8'd12,  9'd113},{  1'b0, 1'b0,   8'd7,   9'd13},{  1'b0, 1'b1,   8'd1,  9'd160}
};
localparam bit [18 : 0] cLARGE_HS_V_TAB_3BY4_PACKED[cLARGE_HS_TAB_3BY4_PACKED_SIZE] = '{
{8'd179, 1'b0,   10'd0},{8'd179, 1'b1, 10'd616},
{8'd178, 1'b0, 10'd602},{8'd178, 1'b1, 10'd617},
{8'd177, 1'b0, 10'd588},{8'd177, 1'b1, 10'd603},
{8'd176, 1'b0, 10'd574},{8'd176, 1'b1, 10'd589},
{8'd175, 1'b0, 10'd560},{8'd175, 1'b1, 10'd575},
{8'd174, 1'b0, 10'd546},{8'd174, 1'b1, 10'd561},
{8'd173, 1'b0, 10'd532},{8'd173, 1'b1, 10'd547},
{8'd172, 1'b0, 10'd518},{8'd172, 1'b1, 10'd533},
{8'd171, 1'b0, 10'd504},{8'd171, 1'b1, 10'd519},
{8'd170, 1'b0, 10'd490},{8'd170, 1'b1, 10'd505},
{8'd169, 1'b0, 10'd476},{8'd169, 1'b1, 10'd491},
{8'd168, 1'b0, 10'd462},{8'd168, 1'b1, 10'd477},
{8'd167, 1'b0, 10'd448},{8'd167, 1'b1, 10'd463},
{8'd166, 1'b0, 10'd434},{8'd166, 1'b1, 10'd449},
{8'd165, 1'b0, 10'd420},{8'd165, 1'b1, 10'd435},
{8'd164, 1'b0, 10'd406},{8'd164, 1'b1, 10'd421},
{8'd163, 1'b0, 10'd392},{8'd163, 1'b1, 10'd407},
{8'd162, 1'b0, 10'd378},{8'd162, 1'b1, 10'd393},
{8'd161, 1'b0, 10'd364},{8'd161, 1'b1, 10'd379},
{8'd160, 1'b0, 10'd350},{8'd160, 1'b1, 10'd365},
{8'd159, 1'b0, 10'd336},{8'd159, 1'b1, 10'd351},
{8'd158, 1'b0, 10'd322},{8'd158, 1'b1, 10'd337},
{8'd157, 1'b0, 10'd308},{8'd157, 1'b1, 10'd323},
{8'd156, 1'b0, 10'd294},{8'd156, 1'b1, 10'd309},
{8'd155, 1'b0, 10'd280},{8'd155, 1'b1, 10'd295},
{8'd154, 1'b0, 10'd266},{8'd154, 1'b1, 10'd281},
{8'd153, 1'b0, 10'd252},{8'd153, 1'b1, 10'd267},
{8'd152, 1'b0, 10'd238},{8'd152, 1'b1, 10'd253},
{8'd151, 1'b0, 10'd224},{8'd151, 1'b1, 10'd239},
{8'd150, 1'b0, 10'd210},{8'd150, 1'b1, 10'd225},
{8'd149, 1'b0, 10'd196},{8'd149, 1'b1, 10'd211},
{8'd148, 1'b0, 10'd182},{8'd148, 1'b1, 10'd197},
{8'd147, 1'b0, 10'd168},{8'd147, 1'b1, 10'd183},
{8'd146, 1'b0, 10'd154},{8'd146, 1'b1, 10'd169},
{8'd145, 1'b0, 10'd140},{8'd145, 1'b1, 10'd155},
{8'd144, 1'b0, 10'd126},{8'd144, 1'b1, 10'd141},
{8'd143, 1'b0, 10'd112},{8'd143, 1'b1, 10'd127},
{8'd142, 1'b0,  10'd98},{8'd142, 1'b1, 10'd113},
{8'd141, 1'b0,  10'd84},{8'd141, 1'b1,  10'd99},
{8'd140, 1'b0,  10'd70},{8'd140, 1'b1,  10'd85},
{8'd139, 1'b0,  10'd56},{8'd139, 1'b1,  10'd71},
{8'd138, 1'b0,  10'd42},{8'd138, 1'b1,  10'd57},
{8'd137, 1'b0,  10'd28},{8'd137, 1'b1,  10'd43},
{8'd136, 1'b0,  10'd14},{8'd136, 1'b1,  10'd29},
{8'd135, 1'b0,   10'd1},{8'd135, 1'b1,  10'd15},
{8'd134, 1'b0,  10'd44},{8'd134, 1'b0, 10'd436},{8'd134, 1'b1, 10'd618},
{8'd133, 1'b0, 10'd338},{8'd133, 1'b0, 10'd520},{8'd133, 1'b1, 10'd604},
{8'd132, 1'b0, 10'd282},{8'd132, 1'b0, 10'd576},{8'd132, 1'b1, 10'd590},
{8'd131, 1'b0,  10'd72},{8'd131, 1'b0, 10'd577},{8'd131, 1'b1, 10'd619},
{8'd130, 1'b0, 10'd464},{8'd130, 1'b0, 10'd534},{8'd130, 1'b1, 10'd562},
{8'd129, 1'b0,  10'd16},{8'd129, 1'b0, 10'd240},{8'd129, 1'b1, 10'd548},
{8'd128, 1'b0, 10'd366},{8'd128, 1'b0, 10'd394},{8'd128, 1'b1, 10'd535},
{8'd127, 1'b0, 10'd268},{8'd127, 1'b0, 10'd450},{8'd127, 1'b1, 10'd521},
{8'd126, 1'b0,   10'd2},{8'd126, 1'b0, 10'd422},{8'd126, 1'b1, 10'd506},
{8'd125, 1'b0, 10'd212},{8'd125, 1'b0, 10'd492},{8'd125, 1'b1, 10'd536},
{8'd124, 1'b0, 10'd339},{8'd124, 1'b0, 10'd478},{8'd124, 1'b1, 10'd507},
{8'd123, 1'b0,  10'd45},{8'd123, 1'b0, 10'd100},{8'd123, 1'b1, 10'd465},
{8'd122, 1'b0, 10'd156},{8'd122, 1'b0, 10'd451},{8'd122, 1'b1, 10'd493},
{8'd121, 1'b0, 10'd254},{8'd121, 1'b0, 10'd437},{8'd121, 1'b1, 10'd563},
{8'd120, 1'b0, 10'd310},{8'd120, 1'b0, 10'd367},{8'd120, 1'b1, 10'd423},
{8'd119, 1'b0, 10'd255},{8'd119, 1'b0, 10'd408},{8'd119, 1'b1, 10'd452},
{8'd118, 1'b0, 10'd352},{8'd118, 1'b0, 10'd380},{8'd118, 1'b1, 10'd395},
{8'd117, 1'b0, 10'd381},{8'd117, 1'b0, 10'd508},{8'd117, 1'b1, 10'd591},
{8'd116, 1'b0, 10'd114},{8'd116, 1'b0, 10'd198},{8'd116, 1'b1, 10'd368},
{8'd115, 1'b0, 10'd353},{8'd115, 1'b0, 10'd605},{8'd115, 1'b1, 10'd606},
{8'd114, 1'b0,  10'd30},{8'd114, 1'b0, 10'd226},{8'd114, 1'b1, 10'd340},
{8'd113, 1'b0,  10'd17},{8'd113, 1'b0, 10'd283},{8'd113, 1'b1, 10'd324},
{8'd112, 1'b0, 10'd311},{8'd112, 1'b0, 10'd396},{8'd112, 1'b1, 10'd494},
{8'd111, 1'b0, 10'd128},{8'd111, 1'b0, 10'd296},{8'd111, 1'b1, 10'd549},
{8'd110, 1'b0, 10'd184},{8'd110, 1'b0, 10'd284},{8'd110, 1'b1, 10'd297},
{8'd109, 1'b0, 10'd269},{8'd109, 1'b0, 10'd325},{8'd109, 1'b1, 10'd479},
{8'd108, 1'b0, 10'd101},{8'd108, 1'b0, 10'd129},{8'd108, 1'b1, 10'd256},
{8'd107, 1'b0,  10'd58},{8'd107, 1'b0, 10'd185},{8'd107, 1'b1, 10'd241},
{8'd106, 1'b0,  10'd86},{8'd106, 1'b0, 10'd227},{8'd106, 1'b1, 10'd326},
{8'd105, 1'b0, 10'd199},{8'd105, 1'b0, 10'd213},{8'd105, 1'b1, 10'd480},
{8'd104, 1'b0, 10'd170},{8'd104, 1'b0, 10'd200},{8'd104, 1'b1, 10'd409},
{8'd103, 1'b0, 10'd186},{8'd103, 1'b0, 10'd298},{8'd103, 1'b1, 10'd564},
{8'd102, 1'b0, 10'd171},{8'd102, 1'b0, 10'd214},{8'd102, 1'b1, 10'd242},
{8'd101, 1'b0, 10'd157},{8'd101, 1'b0, 10'd522},{8'd101, 1'b1, 10'd550},
{8'd100, 1'b0,  10'd59},{8'd100, 1'b0, 10'd142},{8'd100, 1'b1, 10'd143},
{ 8'd99, 1'b0, 10'd130},{ 8'd99, 1'b0, 10'd144},{ 8'd99, 1'b1, 10'd438},
{ 8'd98, 1'b0,  10'd87},{ 8'd98, 1'b0, 10'd115},{ 8'd98, 1'b1, 10'd312},
{ 8'd97, 1'b0, 10'd102},{ 8'd97, 1'b0, 10'd158},{ 8'd97, 1'b1, 10'd382},
{ 8'd96, 1'b0,  10'd88},{ 8'd96, 1'b0, 10'd116},{ 8'd96, 1'b1, 10'd270},
{ 8'd95, 1'b0,  10'd73},{ 8'd95, 1'b0, 10'd466},{ 8'd95, 1'b1, 10'd578},
{ 8'd94, 1'b0,   10'd3},{ 8'd94, 1'b0,  10'd60},{ 8'd94, 1'b1,  10'd74},
{ 8'd93, 1'b0,  10'd46},{ 8'd93, 1'b0, 10'd592},{ 8'd93, 1'b1, 10'd620},
{ 8'd92, 1'b0,  10'd31},{ 8'd92, 1'b0, 10'd354},{ 8'd92, 1'b1, 10'd410},
{ 8'd91, 1'b0,  10'd18},{ 8'd91, 1'b0, 10'd228},{ 8'd91, 1'b1, 10'd424},
{ 8'd90, 1'b0,   10'd4},{ 8'd90, 1'b0,  10'd32},{ 8'd90, 1'b1, 10'd172},
{ 8'd89, 1'b0,  10'd89},{ 8'd89, 1'b0, 10'd117},{ 8'd89, 1'b1, 10'd621},
{ 8'd88, 1'b0, 10'd243},{ 8'd88, 1'b0, 10'd537},{ 8'd88, 1'b1, 10'd607},
{ 8'd87, 1'b0, 10'd131},{ 8'd87, 1'b0, 10'd271},{ 8'd87, 1'b1, 10'd593},
{ 8'd86, 1'b0, 10'd215},{ 8'd86, 1'b0, 10'd495},{ 8'd86, 1'b1, 10'd579},
{ 8'd85, 1'b0,  10'd33},{ 8'd85, 1'b0, 10'd229},{ 8'd85, 1'b1, 10'd565},
{ 8'd84, 1'b0, 10'd230},{ 8'd84, 1'b0, 10'd313},{ 8'd84, 1'b1, 10'd551},
{ 8'd83, 1'b0, 10'd538},{ 8'd83, 1'b0, 10'd552},{ 8'd83, 1'b1, 10'd580},
{ 8'd82, 1'b0,  10'd19},{ 8'd82, 1'b0, 10'd299},{ 8'd82, 1'b1, 10'd523},
{ 8'd81, 1'b0, 10'd314},{ 8'd81, 1'b0, 10'd355},{ 8'd81, 1'b1, 10'd509},
{ 8'd80, 1'b0, 10'd341},{ 8'd80, 1'b0, 10'd411},{ 8'd80, 1'b1, 10'd496},
{ 8'd79, 1'b0, 10'd356},{ 8'd79, 1'b0, 10'd481},{ 8'd79, 1'b1, 10'd510},
{ 8'd78, 1'b0, 10'd145},{ 8'd78, 1'b0, 10'd342},{ 8'd78, 1'b1, 10'd467},
{ 8'd77, 1'b0,  10'd75},{ 8'd77, 1'b0, 10'd272},{ 8'd77, 1'b1, 10'd453},
{ 8'd76, 1'b0, 10'd173},{ 8'd76, 1'b0, 10'd439},{ 8'd76, 1'b1, 10'd524},
{ 8'd75, 1'b0, 10'd397},{ 8'd75, 1'b0, 10'd425},{ 8'd75, 1'b1, 10'd622},
{ 8'd74, 1'b0, 10'd285},{ 8'd74, 1'b0, 10'd412},{ 8'd74, 1'b1, 10'd608},
{ 8'd73, 1'b0,  10'd76},{ 8'd73, 1'b0, 10'd383},{ 8'd73, 1'b1, 10'd398},
{ 8'd72, 1'b0, 10'd384},{ 8'd72, 1'b0, 10'd581},{ 8'd72, 1'b1, 10'd609},
{ 8'd71, 1'b0, 10'd369},{ 8'd71, 1'b0, 10'd399},{ 8'd71, 1'b1, 10'd440},
{ 8'd70, 1'b0, 10'd357},{ 8'd70, 1'b0, 10'd426},{ 8'd70, 1'b1, 10'd454},
{ 8'd69, 1'b0,   10'd5},{ 8'd69, 1'b0, 10'd244},{ 8'd69, 1'b1, 10'd343},
{ 8'd68, 1'b0, 10'd187},{ 8'd68, 1'b0, 10'd216},{ 8'd68, 1'b1, 10'd327},
{ 8'd67, 1'b0, 10'd315},{ 8'd67, 1'b0, 10'd370},{ 8'd67, 1'b1, 10'd566},
{ 8'd66, 1'b0, 10'd103},{ 8'd66, 1'b0, 10'd300},{ 8'd66, 1'b1, 10'd511},
{ 8'd65, 1'b0, 10'd286},{ 8'd65, 1'b0, 10'd427},{ 8'd65, 1'b1, 10'd468},
{ 8'd64, 1'b0, 10'd273},{ 8'd64, 1'b0, 10'd328},{ 8'd64, 1'b1, 10'd539},
{ 8'd63, 1'b0, 10'd146},{ 8'd63, 1'b0, 10'd257},{ 8'd63, 1'b1, 10'd594},
{ 8'd62, 1'b0,  10'd20},{ 8'd62, 1'b0, 10'd201},{ 8'd62, 1'b1, 10'd245},
{ 8'd61, 1'b0, 10'd231},{ 8'd61, 1'b0, 10'd482},{ 8'd61, 1'b1, 10'd567},
{ 8'd60, 1'b0, 10'd217},{ 8'd60, 1'b0, 10'd258},{ 8'd60, 1'b1, 10'd623},
{ 8'd59, 1'b0,   10'd6},{ 8'd59, 1'b0, 10'd202},{ 8'd59, 1'b1, 10'd441},
{ 8'd58, 1'b0, 10'd188},{ 8'd58, 1'b0, 10'd371},{ 8'd58, 1'b1, 10'd483},
{ 8'd57, 1'b0, 10'd132},{ 8'd57, 1'b0, 10'd159},{ 8'd57, 1'b1, 10'd174},
{ 8'd56, 1'b0, 10'd160},{ 8'd56, 1'b0, 10'd161},{ 8'd56, 1'b1, 10'd301},
{ 8'd55, 1'b0, 10'd118},{ 8'd55, 1'b0, 10'd147},{ 8'd55, 1'b1, 10'd329},
{ 8'd54, 1'b0, 10'd133},{ 8'd54, 1'b0, 10'd525},{ 8'd54, 1'b1, 10'd595},
{ 8'd53, 1'b0, 10'd119},{ 8'd53, 1'b0, 10'd189},{ 8'd53, 1'b1, 10'd497},
{ 8'd52, 1'b0, 10'd104},{ 8'd52, 1'b0, 10'd175},{ 8'd52, 1'b1, 10'd469},
{ 8'd51, 1'b0,  10'd34},{ 8'd51, 1'b0,  10'd90},{ 8'd51, 1'b1, 10'd203},
{ 8'd50, 1'b0,  10'd47},{ 8'd50, 1'b0,  10'd77},{ 8'd50, 1'b1, 10'd259},
{ 8'd49, 1'b0,  10'd61},{ 8'd49, 1'b0, 10'd413},{ 8'd49, 1'b1, 10'd553},
{ 8'd48, 1'b0,  10'd48},{ 8'd48, 1'b0,  10'd49},{ 8'd48, 1'b1,  10'd91},
{ 8'd47, 1'b0,  10'd35},{ 8'd47, 1'b0, 10'd105},{ 8'd47, 1'b1, 10'd385},
{ 8'd46, 1'b0,  10'd21},{ 8'd46, 1'b0,  10'd62},{ 8'd46, 1'b1, 10'd287},
{ 8'd45, 1'b0,   10'd7},{ 8'd45, 1'b0,  10'd63},{ 8'd45, 1'b1, 10'd455},
{ 8'd44, 1'b0, 10'd442},{ 8'd44, 1'b0, 10'd582},{ 8'd44, 1'b1, 10'd624},
{ 8'd43, 1'b0, 10'd400},{ 8'd43, 1'b0, 10'd610},{ 8'd43, 1'b1, 10'd625},
{ 8'd42, 1'b0, 10'd358},{ 8'd42, 1'b0, 10'd470},{ 8'd42, 1'b1, 10'd596},
{ 8'd41, 1'b0, 10'd190},{ 8'd41, 1'b0, 10'd583},{ 8'd41, 1'b1, 10'd611},
{ 8'd40, 1'b0,  10'd22},{ 8'd40, 1'b0,  10'd36},{ 8'd40, 1'b1, 10'd568},
{ 8'd39, 1'b0,  10'd23},{ 8'd39, 1'b0, 10'd246},{ 8'd39, 1'b1, 10'd554},
{ 8'd38, 1'b0, 10'd288},{ 8'd38, 1'b0, 10'd344},{ 8'd38, 1'b1, 10'd540},
{ 8'd37, 1'b0, 10'd471},{ 8'd37, 1'b0, 10'd484},{ 8'd37, 1'b1, 10'd526},
{ 8'd36, 1'b0,  10'd64},{ 8'd36, 1'b0, 10'd330},{ 8'd36, 1'b1, 10'd512},
{ 8'd35, 1'b0, 10'd232},{ 8'd35, 1'b0, 10'd274},{ 8'd35, 1'b1, 10'd498},
{ 8'd34, 1'b0, 10'd386},{ 8'd34, 1'b0, 10'd485},{ 8'd34, 1'b1, 10'd486},
{ 8'd33, 1'b0, 10'd106},{ 8'd33, 1'b0, 10'd472},{ 8'd33, 1'b1, 10'd541},
{ 8'd32, 1'b0,  10'd78},{ 8'd32, 1'b0, 10'd456},{ 8'd32, 1'b1, 10'd555},
{ 8'd31, 1'b0,   10'd8},{ 8'd31, 1'b0, 10'd176},{ 8'd31, 1'b1, 10'd443},
{ 8'd30, 1'b0,  10'd37},{ 8'd30, 1'b0,  10'd79},{ 8'd30, 1'b1, 10'd428},
{ 8'd29, 1'b0,  10'd65},{ 8'd29, 1'b0, 10'd134},{ 8'd29, 1'b1, 10'd414},
{ 8'd28, 1'b0, 10'd247},{ 8'd28, 1'b0, 10'd401},{ 8'd28, 1'b1, 10'd513},
{ 8'd27, 1'b0, 10'd289},{ 8'd27, 1'b0, 10'd345},{ 8'd27, 1'b1, 10'd387},
{ 8'd26, 1'b0, 10'd218},{ 8'd26, 1'b0, 10'd372},{ 8'd26, 1'b1, 10'd499},
{ 8'd25, 1'b0, 10'd359},{ 8'd25, 1'b0, 10'd373},{ 8'd25, 1'b1, 10'd402},
{ 8'd24, 1'b0, 10'd346},{ 8'd24, 1'b0, 10'd597},{ 8'd24, 1'b1, 10'd598},
{ 8'd23, 1'b0, 10'd162},{ 8'd23, 1'b0, 10'd331},{ 8'd23, 1'b1, 10'd332},
{ 8'd22, 1'b0, 10'd204},{ 8'd22, 1'b0, 10'd316},{ 8'd22, 1'b1, 10'd360},
{ 8'd21, 1'b0, 10'd120},{ 8'd21, 1'b0, 10'd302},{ 8'd21, 1'b1, 10'd542},
{ 8'd20, 1'b0, 10'd290},{ 8'd20, 1'b0, 10'd388},{ 8'd20, 1'b1, 10'd429},
{ 8'd19, 1'b0, 10'd107},{ 8'd19, 1'b0, 10'd275},{ 8'd19, 1'b1, 10'd556},
{ 8'd18, 1'b0, 10'd219},{ 8'd18, 1'b0, 10'd260},{ 8'd18, 1'b1, 10'd415},
{ 8'd17, 1'b0,  10'd50},{ 8'd17, 1'b0, 10'd248},{ 8'd17, 1'b1, 10'd457},
{ 8'd16, 1'b0,  10'd92},{ 8'd16, 1'b0, 10'd233},{ 8'd16, 1'b1, 10'd303},
{ 8'd15, 1'b0, 10'd163},{ 8'd15, 1'b0, 10'd220},{ 8'd15, 1'b1, 10'd626},
{ 8'd14, 1'b0, 10'd108},{ 8'd14, 1'b0, 10'd205},{ 8'd14, 1'b0, 10'd261},{ 8'd14, 1'b0, 10'd374},{ 8'd14, 1'b0, 10'd375},{ 8'd14, 1'b0, 10'd403},{ 8'd14, 1'b0, 10'd404},{ 8'd14, 1'b0, 10'd473},{ 8'd14, 1'b0, 10'd474},{ 8'd14, 1'b0, 10'd500},{ 8'd14, 1'b0, 10'd527},{ 8'd14, 1'b1, 10'd543},
{ 8'd13, 1'b0, 10'd109},{ 8'd13, 1'b0, 10'd148},{ 8'd13, 1'b0, 10'd177},{ 8'd13, 1'b0, 10'd191},{ 8'd13, 1'b0, 10'd192},{ 8'd13, 1'b0, 10'd206},{ 8'd13, 1'b0, 10'd276},{ 8'd13, 1'b0, 10'd444},{ 8'd13, 1'b0, 10'd514},{ 8'd13, 1'b0, 10'd528},{ 8'd13, 1'b0, 10'd569},{ 8'd13, 1'b1, 10'd584},
{ 8'd12, 1'b0,  10'd93},{ 8'd12, 1'b0, 10'd121},{ 8'd12, 1'b0, 10'd149},{ 8'd12, 1'b0, 10'd178},{ 8'd12, 1'b0, 10'd179},{ 8'd12, 1'b0, 10'd207},{ 8'd12, 1'b0, 10'd277},{ 8'd12, 1'b0, 10'd416},{ 8'd12, 1'b0, 10'd487},{ 8'd12, 1'b0, 10'd529},{ 8'd12, 1'b0, 10'd570},{ 8'd12, 1'b1, 10'd627},
{ 8'd11, 1'b0,  10'd66},{ 8'd11, 1'b0, 10'd164},{ 8'd11, 1'b0, 10'd193},{ 8'd11, 1'b0, 10'd262},{ 8'd11, 1'b0, 10'd304},{ 8'd11, 1'b0, 10'd347},{ 8'd11, 1'b0, 10'd361},{ 8'd11, 1'b0, 10'd417},{ 8'd11, 1'b0, 10'd501},{ 8'd11, 1'b0, 10'd571},{ 8'd11, 1'b0, 10'd585},{ 8'd11, 1'b1, 10'd612},
{ 8'd10, 1'b0,   10'd9},{ 8'd10, 1'b0,  10'd67},{ 8'd10, 1'b0, 10'd122},{ 8'd10, 1'b0, 10'd150},{ 8'd10, 1'b0, 10'd194},{ 8'd10, 1'b0, 10'd221},{ 8'd10, 1'b0, 10'd291},{ 8'd10, 1'b0, 10'd405},{ 8'd10, 1'b0, 10'd430},{ 8'd10, 1'b0, 10'd475},{ 8'd10, 1'b0, 10'd544},{ 8'd10, 1'b1, 10'd557},
{  8'd9, 1'b0,  10'd24},{  8'd9, 1'b0,  10'd80},{  8'd9, 1'b0,  10'd94},{  8'd9, 1'b0, 10'd110},{  8'd9, 1'b0, 10'd135},{  8'd9, 1'b0, 10'd151},{  8'd9, 1'b0, 10'd234},{  8'd9, 1'b0, 10'd317},{  8'd9, 1'b0, 10'd348},{  8'd9, 1'b0, 10'd362},{  8'd9, 1'b0, 10'd389},{  8'd9, 1'b1, 10'd530},
{  8'd8, 1'b0,  10'd51},{  8'd8, 1'b0,  10'd52},{  8'd8, 1'b0,  10'd95},{  8'd8, 1'b0, 10'd123},{  8'd8, 1'b0, 10'd124},{  8'd8, 1'b0, 10'd165},{  8'd8, 1'b0, 10'd292},{  8'd8, 1'b0, 10'd318},{  8'd8, 1'b0, 10'd363},{  8'd8, 1'b0, 10'd390},{  8'd8, 1'b0, 10'd458},{  8'd8, 1'b1, 10'd586},
{  8'd7, 1'b0,  10'd25},{  8'd7, 1'b0,  10'd38},{  8'd7, 1'b0,  10'd53},{  8'd7, 1'b0, 10'd111},{  8'd7, 1'b0, 10'd222},{  8'd7, 1'b0, 10'd263},{  8'd7, 1'b0, 10'd376},{  8'd7, 1'b0, 10'd445},{  8'd7, 1'b0, 10'd488},{  8'd7, 1'b0, 10'd545},{  8'd7, 1'b0, 10'd558},{  8'd7, 1'b1, 10'd628},
{  8'd6, 1'b0,  10'd10},{  8'd6, 1'b0,  10'd96},{  8'd6, 1'b0, 10'd136},{  8'd6, 1'b0, 10'd235},{  8'd6, 1'b0, 10'd236},{  8'd6, 1'b0, 10'd264},{  8'd6, 1'b0, 10'd265},{  8'd6, 1'b0, 10'd333},{  8'd6, 1'b0, 10'd391},{  8'd6, 1'b0, 10'd431},{  8'd6, 1'b0, 10'd432},{  8'd6, 1'b1, 10'd515},
{  8'd5, 1'b0,  10'd54},{  8'd5, 1'b0,  10'd81},{  8'd5, 1'b0,  10'd82},{  8'd5, 1'b0,  10'd83},{  8'd5, 1'b0,  10'd97},{  8'd5, 1'b0, 10'd166},{  8'd5, 1'b0, 10'd293},{  8'd5, 1'b0, 10'd334},{  8'd5, 1'b0, 10'd418},{  8'd5, 1'b0, 10'd502},{  8'd5, 1'b0, 10'd516},{  8'd5, 1'b1, 10'd587},
{  8'd4, 1'b0,  10'd68},{  8'd4, 1'b0, 10'd125},{  8'd4, 1'b0, 10'd137},{  8'd4, 1'b0, 10'd152},{  8'd4, 1'b0, 10'd195},{  8'd4, 1'b0, 10'd208},{  8'd4, 1'b0, 10'd223},{  8'd4, 1'b0, 10'd278},{  8'd4, 1'b0, 10'd305},{  8'd4, 1'b0, 10'd319},{  8'd4, 1'b0, 10'd446},{  8'd4, 1'b1, 10'd613},
{  8'd3, 1'b0,  10'd11},{  8'd3, 1'b0,  10'd26},{  8'd3, 1'b0,  10'd55},{  8'd3, 1'b0, 10'd209},{  8'd3, 1'b0, 10'd237},{  8'd3, 1'b0, 10'd249},{  8'd3, 1'b0, 10'd250},{  8'd3, 1'b0, 10'd433},{  8'd3, 1'b0, 10'd459},{  8'd3, 1'b0, 10'd503},{  8'd3, 1'b0, 10'd517},{  8'd3, 1'b1, 10'd599},
{  8'd2, 1'b0,  10'd12},{  8'd2, 1'b0,  10'd39},{  8'd2, 1'b0,  10'd40},{  8'd2, 1'b0,  10'd69},{  8'd2, 1'b0, 10'd138},{  8'd2, 1'b0, 10'd180},{  8'd2, 1'b0, 10'd251},{  8'd2, 1'b0, 10'd306},{  8'd2, 1'b0, 10'd320},{  8'd2, 1'b0, 10'd460},{  8'd2, 1'b0, 10'd489},{  8'd2, 1'b1, 10'd614},
{  8'd1, 1'b0,  10'd27},{  8'd1, 1'b0,  10'd41},{  8'd1, 1'b0, 10'd139},{  8'd1, 1'b0, 10'd153},{  8'd1, 1'b0, 10'd279},{  8'd1, 1'b0, 10'd307},{  8'd1, 1'b0, 10'd461},{  8'd1, 1'b0, 10'd531},{  8'd1, 1'b0, 10'd600},{  8'd1, 1'b0, 10'd601},{  8'd1, 1'b0, 10'd615},{  8'd1, 1'b1, 10'd629},
{  8'd0, 1'b0,  10'd13},{  8'd0, 1'b0, 10'd167},{  8'd0, 1'b0, 10'd181},{  8'd0, 1'b0, 10'd321},{  8'd0, 1'b0, 10'd335},{  8'd0, 1'b0, 10'd349},{  8'd0, 1'b0, 10'd377},{  8'd0, 1'b0, 10'd419},{  8'd0, 1'b0, 10'd447},{  8'd0, 1'b0, 10'd559},{  8'd0, 1'b0, 10'd572},{  8'd0, 1'b1, 10'd573}
};
localparam int          cLARGE_HS_TAB_4BY5_PACKED_SIZE = 648;
localparam bit [18 : 0] cLARGE_HS_TAB_4BY5_PACKED[cLARGE_HS_TAB_4BY5_PACKED_SIZE] = '{
{  1'b1, 1'b0, 8'd179,    9'd1},{  1'b0, 1'b0, 8'd144,    9'd0},{  1'b0, 1'b0, 8'd139,  9'd258},{  1'b0, 1'b0, 8'd125,  9'd231},{  1'b0, 1'b0, 8'd108,    9'd0},{  1'b0, 1'b0,  8'd86,  9'd200},{  1'b0, 1'b0,  8'd81,   9'd34},{  1'b0, 1'b0,  8'd72,    9'd0},{  1'b0, 1'b0,  8'd49,   9'd72},{  1'b0, 1'b0,  8'd39,   9'd61},{  1'b0, 1'b0,  8'd36,    9'd0},{  1'b0, 1'b0,  8'd25,  9'd121},{  1'b0, 1'b0,  8'd17,  9'd243},{  1'b0, 1'b0,  8'd15,  9'd319},{  1'b0, 1'b0,  8'd15,  9'd181},{  1'b0, 1'b0,  8'd12,  9'd325},{  1'b0, 1'b0,   8'd6,  9'd104},{  1'b0, 1'b1,   8'd0,    9'd0},
{  1'b0, 1'b0, 8'd145,    9'd0},{  1'b0, 1'b0, 8'd144,    9'd0},{  1'b0, 1'b0, 8'd121,  9'd211},{  1'b0, 1'b0, 8'd118,  9'd344},{  1'b0, 1'b0, 8'd109,    9'd0},{  1'b0, 1'b0,  8'd98,  9'd359},{  1'b0, 1'b0,  8'd96,   9'd23},{  1'b0, 1'b0,  8'd73,    9'd0},{  1'b0, 1'b0,  8'd63,   9'd97},{  1'b0, 1'b0,  8'd41,  9'd297},{  1'b0, 1'b0,  8'd37,    9'd0},{  1'b0, 1'b0,  8'd33,  9'd289},{  1'b0, 1'b0,  8'd27,  9'd330},{  1'b0, 1'b0,  8'd17,  9'd315},{  1'b0, 1'b0,  8'd14,   9'd96},{  1'b0, 1'b0,  8'd10,  9'd242},{  1'b0, 1'b0,   8'd9,    9'd7},{  1'b0, 1'b1,   8'd1,    9'd0},
{  1'b0, 1'b0, 8'd146,    9'd0},{  1'b0, 1'b0, 8'd145,    9'd0},{  1'b0, 1'b0, 8'd125,  9'd183},{  1'b0, 1'b0, 8'd118,  9'd333},{  1'b0, 1'b0, 8'd110,    9'd0},{  1'b0, 1'b0, 8'd106,  9'd226},{  1'b0, 1'b0,  8'd78,  9'd156},{  1'b0, 1'b0,  8'd74,    9'd0},{  1'b0, 1'b0,  8'd67,   9'd58},{  1'b0, 1'b0,  8'd48,  9'd332},{  1'b0, 1'b0,  8'd38,    9'd0},{  1'b0, 1'b0,  8'd21,  9'd341},{  1'b0, 1'b0,  8'd19,   9'd28},{  1'b0, 1'b0,  8'd12,  9'd107},{  1'b0, 1'b0,  8'd10,  9'd218},{  1'b0, 1'b0,   8'd7,   9'd31},{  1'b0, 1'b0,   8'd5,   9'd95},{  1'b0, 1'b1,   8'd2,    9'd0},
{  1'b0, 1'b0, 8'd147,    9'd0},{  1'b0, 1'b0, 8'd146,    9'd0},{  1'b0, 1'b0, 8'd129,  9'd162},{  1'b0, 1'b0, 8'd128,    9'd7},{  1'b0, 1'b0, 8'd111,    9'd0},{  1'b0, 1'b0,  8'd94,  9'd184},{  1'b0, 1'b0,  8'd75,    9'd0},{  1'b0, 1'b0,  8'd72,  9'd137},{  1'b0, 1'b0,  8'd58,  9'd216},{  1'b0, 1'b0,  8'd40,  9'd209},{  1'b0, 1'b0,  8'd39,    9'd0},{  1'b0, 1'b0,  8'd18,  9'd282},{  1'b0, 1'b0,  8'd15,   9'd76},{  1'b0, 1'b0,  8'd11,  9'd254},{  1'b0, 1'b0,   8'd9,   9'd65},{  1'b0, 1'b0,   8'd5,   9'd59},{  1'b0, 1'b0,   8'd5,   9'd28},{  1'b0, 1'b1,   8'd3,    9'd0},
{  1'b0, 1'b0, 8'd148,    9'd0},{  1'b0, 1'b0, 8'd147,    9'd0},{  1'b0, 1'b0, 8'd134,  9'd270},{  1'b0, 1'b0, 8'd122,    9'd3},{  1'b0, 1'b0, 8'd112,    9'd0},{  1'b0, 1'b0, 8'd104,   9'd17},{  1'b0, 1'b0,  8'd84,   9'd90},{  1'b0, 1'b0,  8'd76,    9'd0},{  1'b0, 1'b0,  8'd54,  9'd167},{  1'b0, 1'b0,  8'd49,  9'd206},{  1'b0, 1'b0,  8'd40,    9'd0},{  1'b0, 1'b0,  8'd31,  9'd176},{  1'b0, 1'b0,  8'd30,   9'd62},{  1'b0, 1'b0,  8'd15,  9'd184},{  1'b0, 1'b0,   8'd7,  9'd180},{  1'b0, 1'b0,   8'd6,   9'd26},{  1'b0, 1'b0,   8'd4,    9'd0},{  1'b0, 1'b1,   8'd4,  9'd333},
{  1'b0, 1'b0, 8'd149,    9'd0},{  1'b0, 1'b0, 8'd148,    9'd0},{  1'b0, 1'b0, 8'd129,  9'd172},{  1'b0, 1'b0, 8'd128,    9'd3},{  1'b0, 1'b0, 8'd113,    9'd0},{  1'b0, 1'b0, 8'd105,  9'd271},{  1'b0, 1'b0,  8'd97,   9'd61},{  1'b0, 1'b0,  8'd77,    9'd0},{  1'b0, 1'b0,  8'd51,   9'd19},{  1'b0, 1'b0,  8'd44,  9'd223},{  1'b0, 1'b0,  8'd41,    9'd0},{  1'b0, 1'b0,  8'd22,  9'd122},{  1'b0, 1'b0,  8'd16,  9'd229},{  1'b0, 1'b0,  8'd13,  9'd318},{  1'b0, 1'b0,   8'd9,  9'd125},{  1'b0, 1'b0,   8'd5,    9'd0},{  1'b0, 1'b0,   8'd5,  9'd113},{  1'b0, 1'b1,   8'd0,    9'd4},
{  1'b0, 1'b0, 8'd150,    9'd0},{  1'b0, 1'b0, 8'd149,    9'd0},{  1'b0, 1'b0, 8'd135,  9'd320},{  1'b0, 1'b0, 8'd132,  9'd152},{  1'b0, 1'b0, 8'd114,    9'd0},{  1'b0, 1'b0,  8'd88,  9'd342},{  1'b0, 1'b0,  8'd88,   9'd61},{  1'b0, 1'b0,  8'd78,    9'd0},{  1'b0, 1'b0,  8'd57,  9'd111},{  1'b0, 1'b0,  8'd42,    9'd0},{  1'b0, 1'b0,  8'd42,   9'd75},{  1'b0, 1'b0,  8'd27,   9'd70},{  1'b0, 1'b0,  8'd13,   9'd69},{  1'b0, 1'b0,  8'd11,   9'd63},{  1'b0, 1'b0,  8'd11,  9'd168},{  1'b0, 1'b0,   8'd8,  9'd234},{  1'b0, 1'b0,   8'd7,  9'd218},{  1'b0, 1'b1,   8'd6,    9'd0},
{  1'b0, 1'b0, 8'd151,    9'd0},{  1'b0, 1'b0, 8'd150,    9'd0},{  1'b0, 1'b0, 8'd136,  9'd264},{  1'b0, 1'b0, 8'd116,  9'd206},{  1'b0, 1'b0, 8'd115,    9'd0},{  1'b0, 1'b0,  8'd86,   9'd91},{  1'b0, 1'b0,  8'd79,    9'd0},{  1'b0, 1'b0,  8'd73,  9'd117},{  1'b0, 1'b0,  8'd63,   9'd68},{  1'b0, 1'b0,  8'd45,  9'd123},{  1'b0, 1'b0,  8'd43,    9'd0},{  1'b0, 1'b0,  8'd19,  9'd291},{  1'b0, 1'b0,  8'd14,  9'd175},{  1'b0, 1'b0,  8'd10,  9'd188},{  1'b0, 1'b0,  8'd10,  9'd227},{  1'b0, 1'b0,   8'd7,    9'd0},{  1'b0, 1'b0,   8'd6,   9'd78},{  1'b0, 1'b1,   8'd4,  9'd335},
{  1'b0, 1'b0, 8'd152,    9'd0},{  1'b0, 1'b0, 8'd151,    9'd0},{  1'b0, 1'b0, 8'd133,   9'd59},{  1'b0, 1'b0, 8'd116,    9'd0},{  1'b0, 1'b0, 8'd112,   9'd96},{  1'b0, 1'b0, 8'd100,  9'd165},{  1'b0, 1'b0,  8'd80,    9'd0},{  1'b0, 1'b0,  8'd77,  9'd249},{  1'b0, 1'b0,  8'd70,  9'd236},{  1'b0, 1'b0,  8'd52,   9'd36},{  1'b0, 1'b0,  8'd44,    9'd0},{  1'b0, 1'b0,  8'd20,  9'd247},{  1'b0, 1'b0,  8'd14,  9'd105},{  1'b0, 1'b0,  8'd10,  9'd248},{  1'b0, 1'b0,   8'd9,   9'd43},{  1'b0, 1'b0,   8'd8,    9'd0},{  1'b0, 1'b0,   8'd8,  9'd262},{  1'b0, 1'b1,   8'd0,  9'd225},
{  1'b0, 1'b0, 8'd153,    9'd0},{  1'b0, 1'b0, 8'd152,    9'd0},{  1'b0, 1'b0, 8'd143,  9'd154},{  1'b0, 1'b0, 8'd123,  9'd221},{  1'b0, 1'b0, 8'd117,    9'd0},{  1'b0, 1'b0, 8'd106,  9'd288},{  1'b0, 1'b0,  8'd99,  9'd243},{  1'b0, 1'b0,  8'd81,    9'd0},{  1'b0, 1'b0,  8'd60,  9'd110},{  1'b0, 1'b0,  8'd45,    9'd0},{  1'b0, 1'b0,  8'd36,  9'd267},{  1'b0, 1'b0,  8'd26,  9'd198},{  1'b0, 1'b0,  8'd13,  9'd162},{  1'b0, 1'b0,   8'd9,    9'd0},{  1'b0, 1'b0,   8'd2,  9'd154},{  1'b0, 1'b0,   8'd2,  9'd291},{  1'b0, 1'b0,   8'd1,  9'd286},{  1'b0, 1'b1,   8'd0,  9'd236},
{  1'b0, 1'b0, 8'd154,    9'd0},{  1'b0, 1'b0, 8'd153,    9'd0},{  1'b0, 1'b0, 8'd122,   9'd40},{  1'b0, 1'b0, 8'd120,  9'd282},{  1'b0, 1'b0, 8'd118,    9'd0},{  1'b0, 1'b0,  8'd92,  9'd286},{  1'b0, 1'b0,  8'd82,    9'd0},{  1'b0, 1'b0,  8'd81,  9'd246},{  1'b0, 1'b0,  8'd65,  9'd183},{  1'b0, 1'b0,  8'd47,  9'd182},{  1'b0, 1'b0,  8'd46,    9'd0},{  1'b0, 1'b0,  8'd25,  9'd264},{  1'b0, 1'b0,  8'd13,  9'd332},{  1'b0, 1'b0,  8'd12,  9'd110},{  1'b0, 1'b0,  8'd12,   9'd60},{  1'b0, 1'b0,  8'd10,    9'd0},{  1'b0, 1'b0,   8'd4,  9'd171},{  1'b0, 1'b1,   8'd3,   9'd90},
{  1'b0, 1'b0, 8'd155,    9'd0},{  1'b0, 1'b0, 8'd154,    9'd0},{  1'b0, 1'b0, 8'd136,  9'd342},{  1'b0, 1'b0, 8'd126,  9'd250},{  1'b0, 1'b0, 8'd119,    9'd0},{  1'b0, 1'b0,  8'd90,  9'd266},{  1'b0, 1'b0,  8'd83,    9'd0},{  1'b0, 1'b0,  8'd75,  9'd151},{  1'b0, 1'b0,  8'd65,  9'd319},{  1'b0, 1'b0,  8'd56,  9'd123},{  1'b0, 1'b0,  8'd47,    9'd0},{  1'b0, 1'b0,  8'd33,  9'd324},{  1'b0, 1'b0,  8'd15,  9'd336},{  1'b0, 1'b0,  8'd15,   9'd15},{  1'b0, 1'b0,  8'd12,  9'd358},{  1'b0, 1'b0,  8'd11,    9'd0},{  1'b0, 1'b0,   8'd8,  9'd114},{  1'b0, 1'b1,   8'd8,  9'd238},
{  1'b0, 1'b0, 8'd156,    9'd0},{  1'b0, 1'b0, 8'd155,    9'd0},{  1'b0, 1'b0, 8'd134,   9'd38},{  1'b0, 1'b0, 8'd120,    9'd0},{  1'b0, 1'b0, 8'd113,  9'd193},{  1'b0, 1'b0,  8'd85,  9'd162},{  1'b0, 1'b0,  8'd84,    9'd0},{  1'b0, 1'b0,  8'd80,  9'd246},{  1'b0, 1'b0,  8'd61,  9'd121},{  1'b0, 1'b0,  8'd48,    9'd0},{  1'b0, 1'b0,  8'd46,  9'd256},{  1'b0, 1'b0,  8'd30,  9'd242},{  1'b0, 1'b0,  8'd12,    9'd0},{  1'b0, 1'b0,  8'd11,  9'd245},{  1'b0, 1'b0,  8'd10,   9'd47},{  1'b0, 1'b0,   8'd2,   9'd78},{  1'b0, 1'b0,   8'd0,   9'd11},{  1'b0, 1'b1,   8'd0,  9'd356},
{  1'b0, 1'b0, 8'd157,    9'd0},{  1'b0, 1'b0, 8'd156,    9'd0},{  1'b0, 1'b0, 8'd131,   9'd97},{  1'b0, 1'b0, 8'd121,    9'd0},{  1'b0, 1'b0, 8'd108,  9'd202},{  1'b0, 1'b0,  8'd85,    9'd0},{  1'b0, 1'b0,  8'd83,  9'd122},{  1'b0, 1'b0,  8'd76,   9'd89},{  1'b0, 1'b0,  8'd70,   9'd51},{  1'b0, 1'b0,  8'd67,  9'd267},{  1'b0, 1'b0,  8'd49,    9'd0},{  1'b0, 1'b0,  8'd29,  9'd303},{  1'b0, 1'b0,  8'd16,   9'd50},{  1'b0, 1'b0,  8'd13,    9'd0},{  1'b0, 1'b0,   8'd9,  9'd157},{  1'b0, 1'b0,   8'd7,  9'd126},{  1'b0, 1'b0,   8'd4,  9'd143},{  1'b0, 1'b1,   8'd3,   9'd14},
{  1'b0, 1'b0, 8'd158,    9'd0},{  1'b0, 1'b0, 8'd157,    9'd0},{  1'b0, 1'b0, 8'd130,  9'd358},{  1'b0, 1'b0, 8'd127,  9'd261},{  1'b0, 1'b0, 8'd122,    9'd0},{  1'b0, 1'b0,  8'd87,  9'd313},{  1'b0, 1'b0,  8'd86,    9'd0},{  1'b0, 1'b0,  8'd83,    9'd7},{  1'b0, 1'b0,  8'd69,   9'd99},{  1'b0, 1'b0,  8'd62,  9'd148},{  1'b0, 1'b0,  8'd50,    9'd0},{  1'b0, 1'b0,  8'd32,  9'd238},{  1'b0, 1'b0,  8'd22,  9'd196},{  1'b0, 1'b0,  8'd17,   9'd58},{  1'b0, 1'b0,  8'd15,  9'd226},{  1'b0, 1'b0,  8'd14,    9'd0},{  1'b0, 1'b0,  8'd11,  9'd331},{  1'b0, 1'b1,   8'd7,   9'd35},
{  1'b0, 1'b0, 8'd159,    9'd0},{  1'b0, 1'b0, 8'd158,    9'd0},{  1'b0, 1'b0, 8'd123,    9'd0},{  1'b0, 1'b0, 8'd121,   9'd37},{  1'b0, 1'b0, 8'd111,  9'd231},{  1'b0, 1'b0, 8'd107,  9'd161},{  1'b0, 1'b0,  8'd99,   9'd59},{  1'b0, 1'b0,  8'd87,    9'd0},{  1'b0, 1'b0,  8'd68,  9'd131},{  1'b0, 1'b0,  8'd57,  9'd265},{  1'b0, 1'b0,  8'd51,    9'd0},{  1'b0, 1'b0,  8'd15,    9'd0},{  1'b0, 1'b0,  8'd12,  9'd203},{  1'b0, 1'b0,  8'd11,  9'd252},{  1'b0, 1'b0,   8'd7,  9'd326},{  1'b0, 1'b0,   8'd7,  9'd112},{  1'b0, 1'b0,   8'd5,  9'd197},{  1'b0, 1'b1,   8'd3,  9'd131},
{  1'b0, 1'b0, 8'd160,    9'd0},{  1'b0, 1'b0, 8'd159,    9'd0},{  1'b0, 1'b0, 8'd143,  9'd197},{  1'b0, 1'b0, 8'd141,    9'd7},{  1'b0, 1'b0, 8'd124,    9'd0},{  1'b0, 1'b0, 8'd100,  9'd333},{  1'b0, 1'b0,  8'd88,    9'd0},{  1'b0, 1'b0,  8'd78,  9'd346},{  1'b0, 1'b0,  8'd69,   9'd72},{  1'b0, 1'b0,  8'd62,  9'd175},{  1'b0, 1'b0,  8'd52,    9'd0},{  1'b0, 1'b0,  8'd17,  9'd186},{  1'b0, 1'b0,  8'd16,    9'd0},{  1'b0, 1'b0,  8'd15,   9'd71},{  1'b0, 1'b0,  8'd11,  9'd325},{  1'b0, 1'b0,   8'd6,  9'd300},{  1'b0, 1'b0,   8'd5,  9'd103},{  1'b0, 1'b1,   8'd0,  9'd311},
{  1'b0, 1'b0, 8'd161,    9'd0},{  1'b0, 1'b0, 8'd160,    9'd0},{  1'b0, 1'b0, 8'd125,    9'd0},{  1'b0, 1'b0, 8'd124,  9'd248},{  1'b0, 1'b0, 8'd124,  9'd205},{  1'b0, 1'b0,  8'd96,  9'd269},{  1'b0, 1'b0,  8'd89,    9'd0},{  1'b0, 1'b0,  8'd79,   9'd40},{  1'b0, 1'b0,  8'd68,   9'd64},{  1'b0, 1'b0,  8'd53,    9'd0},{  1'b0, 1'b0,  8'd46,  9'd115},{  1'b0, 1'b0,  8'd17,    9'd0},{  1'b0, 1'b0,  8'd17,  9'd152},{  1'b0, 1'b0,   8'd8,   9'd11},{  1'b0, 1'b0,   8'd6,  9'd321},{  1'b0, 1'b0,   8'd1,  9'd145},{  1'b0, 1'b0,   8'd1,  9'd107},{  1'b0, 1'b1,   8'd1,   9'd97},
{  1'b0, 1'b0, 8'd162,    9'd0},{  1'b0, 1'b0, 8'd161,    9'd0},{  1'b0, 1'b0, 8'd127,  9'd171},{  1'b0, 1'b0, 8'd126,    9'd0},{  1'b0, 1'b0, 8'd123,  9'd235},{  1'b0, 1'b0, 8'd104,  9'd198},{  1'b0, 1'b0,  8'd93,  9'd307},{  1'b0, 1'b0,  8'd90,    9'd0},{  1'b0, 1'b0,  8'd59,   9'd41},{  1'b0, 1'b0,  8'd54,    9'd0},{  1'b0, 1'b0,  8'd53,  9'd331},{  1'b0, 1'b0,  8'd35,   9'd88},{  1'b0, 1'b0,  8'd18,    9'd0},{  1'b0, 1'b0,  8'd16,  9'd181},{  1'b0, 1'b0,  8'd12,  9'd229},{  1'b0, 1'b0,   8'd9,  9'd253},{  1'b0, 1'b0,   8'd8,  9'd344},{  1'b0, 1'b1,   8'd0,  9'd278},
{  1'b0, 1'b0, 8'd163,    9'd0},{  1'b0, 1'b0, 8'd162,    9'd0},{  1'b0, 1'b0, 8'd127,    9'd0},{  1'b0, 1'b0, 8'd119,  9'd270},{  1'b0, 1'b0, 8'd110,  9'd250},{  1'b0, 1'b0,  8'd97,   9'd50},{  1'b0, 1'b0,  8'd91,    9'd0},{  1'b0, 1'b0,  8'd82,  9'd232},{  1'b0, 1'b0,  8'd55,    9'd0},{  1'b0, 1'b0,  8'd54,  9'd265},{  1'b0, 1'b0,  8'd38,  9'd135},{  1'b0, 1'b0,  8'd21,  9'd284},{  1'b0, 1'b0,  8'd19,    9'd0},{  1'b0, 1'b0,  8'd16,  9'd128},{  1'b0, 1'b0,  8'd11,  9'd151},{  1'b0, 1'b0,   8'd5,  9'd159},{  1'b0, 1'b0,   8'd4,   9'd37},{  1'b0, 1'b1,   8'd2,  9'd216},
{  1'b0, 1'b0, 8'd164,    9'd0},{  1'b0, 1'b0, 8'd163,    9'd0},{  1'b0, 1'b0, 8'd139,   9'd85},{  1'b0, 1'b0, 8'd128,    9'd0},{  1'b0, 1'b0, 8'd117,  9'd225},{  1'b0, 1'b0, 8'd107,  9'd211},{  1'b0, 1'b0,  8'd92,    9'd0},{  1'b0, 1'b0,  8'd79,   9'd35},{  1'b0, 1'b0,  8'd56,    9'd0},{  1'b0, 1'b0,  8'd52,   9'd25},{  1'b0, 1'b0,  8'd39,    9'd9},{  1'b0, 1'b0,  8'd29,   9'd84},{  1'b0, 1'b0,  8'd20,    9'd0},{  1'b0, 1'b0,  8'd17,   9'd81},{  1'b0, 1'b0,  8'd14,  9'd221},{  1'b0, 1'b0,   8'd3,  9'd119},{  1'b0, 1'b0,   8'd2,  9'd336},{  1'b0, 1'b1,   8'd2,   9'd82},
{  1'b0, 1'b0, 8'd165,    9'd0},{  1'b0, 1'b0, 8'd164,    9'd0},{  1'b0, 1'b0, 8'd131,  9'd121},{  1'b0, 1'b0, 8'd129,    9'd0},{  1'b0, 1'b0, 8'd116,  9'd155},{  1'b0, 1'b0,  8'd93,    9'd0},{  1'b0, 1'b0,  8'd92,  9'd334},{  1'b0, 1'b0,  8'd77,   9'd18},{  1'b0, 1'b0,  8'd60,  9'd298},{  1'b0, 1'b0,  8'd57,    9'd0},{  1'b0, 1'b0,  8'd56,  9'd116},{  1'b0, 1'b0,  8'd26,  9'd285},{  1'b0, 1'b0,  8'd21,    9'd0},{  1'b0, 1'b0,  8'd17,  9'd345},{  1'b0, 1'b0,  8'd14,  9'd214},{  1'b0, 1'b0,  8'd14,  9'd166},{  1'b0, 1'b0,  8'd13,  9'd311},{  1'b0, 1'b1,   8'd1,  9'd296},
{  1'b0, 1'b0, 8'd166,    9'd0},{  1'b0, 1'b0, 8'd165,    9'd0},{  1'b0, 1'b0, 8'd138,  9'd250},{  1'b0, 1'b0, 8'd130,    9'd0},{  1'b0, 1'b0, 8'd111,  9'd122},{  1'b0, 1'b0,  8'd94,    9'd0},{  1'b0, 1'b0,  8'd76,  9'd156},{  1'b0, 1'b0,  8'd75,  9'd193},{  1'b0, 1'b0,  8'd58,    9'd0},{  1'b0, 1'b0,  8'd45,  9'd134},{  1'b0, 1'b0,  8'd43,  9'd166},{  1'b0, 1'b0,  8'd22,    9'd0},{  1'b0, 1'b0,  8'd16,  9'd168},{  1'b0, 1'b0,  8'd16,  9'd103},{  1'b0, 1'b0,  8'd16,  9'd329},{  1'b0, 1'b0,   8'd6,  9'd264},{  1'b0, 1'b0,   8'd6,  9'd319},{  1'b0, 1'b1,   8'd1,   9'd13},
{  1'b0, 1'b0, 8'd167,    9'd0},{  1'b0, 1'b0, 8'd166,    9'd0},{  1'b0, 1'b0, 8'd137,  9'd228},{  1'b0, 1'b0, 8'd131,    9'd0},{  1'b0, 1'b0, 8'd113,   9'd56},{  1'b0, 1'b0, 8'd101,   9'd88},{  1'b0, 1'b0,  8'd95,    9'd0},{  1'b0, 1'b0,  8'd89,  9'd125},{  1'b0, 1'b0,  8'd61,   9'd96},{  1'b0, 1'b0,  8'd59,    9'd0},{  1'b0, 1'b0,  8'd42,  9'd187},{  1'b0, 1'b0,  8'd34,  9'd179},{  1'b0, 1'b0,  8'd23,    9'd0},{  1'b0, 1'b0,   8'd7,  9'd319},{  1'b0, 1'b0,   8'd7,  9'd144},{  1'b0, 1'b0,   8'd7,  9'd355},{  1'b0, 1'b0,   8'd4,  9'd338},{  1'b0, 1'b1,   8'd4,   9'd65},
{  1'b0, 1'b0, 8'd168,    9'd0},{  1'b0, 1'b0, 8'd167,    9'd0},{  1'b0, 1'b0, 8'd137,   9'd48},{  1'b0, 1'b0, 8'd132,    9'd0},{  1'b0, 1'b0, 8'd109,  9'd215},{  1'b0, 1'b0, 8'd103,  9'd197},{  1'b0, 1'b0,  8'd96,    9'd0},{  1'b0, 1'b0,  8'd74,  9'd304},{  1'b0, 1'b0,  8'd60,    9'd0},{  1'b0, 1'b0,  8'd55,    9'd8},{  1'b0, 1'b0,  8'd50,  9'd267},{  1'b0, 1'b0,  8'd24,    9'd0},{  1'b0, 1'b0,  8'd15,  9'd273},{  1'b0, 1'b0,  8'd11,  9'd120},{  1'b0, 1'b0,   8'd5,  9'd189},{  1'b0, 1'b0,   8'd5,  9'd306},{  1'b0, 1'b0,   8'd2,   9'd15},{  1'b0, 1'b1,   8'd0,  9'd176},
{  1'b0, 1'b0, 8'd169,    9'd0},{  1'b0, 1'b0, 8'd168,    9'd0},{  1'b0, 1'b0, 8'd133,    9'd0},{  1'b0, 1'b0, 8'd133,  9'd123},{  1'b0, 1'b0, 8'd117,  9'd135},{  1'b0, 1'b0, 8'd102,  9'd303},{  1'b0, 1'b0,  8'd97,    9'd0},{  1'b0, 1'b0,  8'd95,  9'd274},{  1'b0, 1'b0,  8'd64,  9'd337},{  1'b0, 1'b0,  8'd64,  9'd205},{  1'b0, 1'b0,  8'd61,    9'd0},{  1'b0, 1'b0,  8'd28,   9'd54},{  1'b0, 1'b0,  8'd25,    9'd0},{  1'b0, 1'b0,  8'd17,  9'd217},{  1'b0, 1'b0,  8'd17,  9'd332},{  1'b0, 1'b0,  8'd14,  9'd125},{  1'b0, 1'b0,  8'd13,   9'd22},{  1'b0, 1'b1,   8'd3,  9'd280},
{  1'b0, 1'b0, 8'd170,    9'd0},{  1'b0, 1'b0, 8'd169,    9'd0},{  1'b0, 1'b0, 8'd134,    9'd0},{  1'b0, 1'b0, 8'd119,  9'd278},{  1'b0, 1'b0, 8'd115,   9'd19},{  1'b0, 1'b0,  8'd98,    9'd0},{  1'b0, 1'b0,  8'd87,   9'd41},{  1'b0, 1'b0,  8'd74,  9'd223},{  1'b0, 1'b0,  8'd62,    9'd0},{  1'b0, 1'b0,  8'd50,  9'd244},{  1'b0, 1'b0,  8'd40,  9'd184},{  1'b0, 1'b0,  8'd26,    9'd0},{  1'b0, 1'b0,  8'd20,  9'd284},{  1'b0, 1'b0,  8'd13,  9'd122},{  1'b0, 1'b0,  8'd10,  9'd228},{  1'b0, 1'b0,   8'd9,  9'd115},{  1'b0, 1'b0,   8'd6,   9'd40},{  1'b0, 1'b1,   8'd1,  9'd103},
{  1'b0, 1'b0, 8'd171,    9'd0},{  1'b0, 1'b0, 8'd170,    9'd0},{  1'b0, 1'b0, 8'd142,  9'd111},{  1'b0, 1'b0, 8'd140,  9'd208},{  1'b0, 1'b0, 8'd135,    9'd0},{  1'b0, 1'b0,  8'd99,    9'd0},{  1'b0, 1'b0,  8'd90,  9'd194},{  1'b0, 1'b0,  8'd85,  9'd167},{  1'b0, 1'b0,  8'd66,  9'd123},{  1'b0, 1'b0,  8'd63,    9'd0},{  1'b0, 1'b0,  8'd44,  9'd306},{  1'b0, 1'b0,  8'd27,    9'd0},{  1'b0, 1'b0,  8'd15,  9'd111},{  1'b0, 1'b0,  8'd13,   9'd40},{  1'b0, 1'b0,  8'd10,  9'd246},{  1'b0, 1'b0,   8'd9,  9'd130},{  1'b0, 1'b0,   8'd8,  9'd123},{  1'b0, 1'b1,   8'd6,  9'd312},
{  1'b0, 1'b0, 8'd172,    9'd0},{  1'b0, 1'b0, 8'd171,    9'd0},{  1'b0, 1'b0, 8'd136,    9'd0},{  1'b0, 1'b0, 8'd130,  9'd106},{  1'b0, 1'b0, 8'd120,   9'd11},{  1'b0, 1'b0, 8'd101,  9'd241},{  1'b0, 1'b0, 8'd100,    9'd0},{  1'b0, 1'b0,  8'd93,  9'd141},{  1'b0, 1'b0,  8'd64,    9'd0},{  1'b0, 1'b0,  8'd58,  9'd339},{  1'b0, 1'b0,  8'd41,   9'd67},{  1'b0, 1'b0,  8'd28,    9'd0},{  1'b0, 1'b0,  8'd24,  9'd332},{  1'b0, 1'b0,  8'd17,  9'd212},{  1'b0, 1'b0,   8'd6,   9'd33},{  1'b0, 1'b0,   8'd5,  9'd298},{  1'b0, 1'b0,   8'd3,   9'd19},{  1'b0, 1'b1,   8'd3,  9'd208},
{  1'b0, 1'b0, 8'd173,    9'd0},{  1'b0, 1'b0, 8'd172,    9'd0},{  1'b0, 1'b0, 8'd142,  9'd342},{  1'b0, 1'b0, 8'd138,   9'd13},{  1'b0, 1'b0, 8'd137,    9'd0},{  1'b0, 1'b0, 8'd101,    9'd0},{  1'b0, 1'b0,  8'd98,  9'd185},{  1'b0, 1'b0,  8'd89,   9'd26},{  1'b0, 1'b0,  8'd65,    9'd0},{  1'b0, 1'b0,  8'd55,  9'd210},{  1'b0, 1'b0,  8'd53,   9'd34},{  1'b0, 1'b0,  8'd29,    9'd0},{  1'b0, 1'b0,  8'd28,  9'd318},{  1'b0, 1'b0,  8'd16,  9'd219},{  1'b0, 1'b0,  8'd14,   9'd42},{  1'b0, 1'b0,  8'd13,   9'd14},{  1'b0, 1'b0,  8'd12,  9'd263},{  1'b0, 1'b1,   8'd2,  9'd196},
{  1'b0, 1'b0, 8'd174,    9'd0},{  1'b0, 1'b0, 8'd173,    9'd0},{  1'b0, 1'b0, 8'd138,    9'd0},{  1'b0, 1'b0, 8'd114,   9'd21},{  1'b0, 1'b0, 8'd112,   9'd17},{  1'b0, 1'b0, 8'd105,  9'd142},{  1'b0, 1'b0, 8'd102,    9'd0},{  1'b0, 1'b0,  8'd94,  9'd191},{  1'b0, 1'b0,  8'd66,    9'd0},{  1'b0, 1'b0,  8'd51,  9'd150},{  1'b0, 1'b0,  8'd47,  9'd340},{  1'b0, 1'b0,  8'd35,  9'd338},{  1'b0, 1'b0,  8'd30,    9'd0},{  1'b0, 1'b0,  8'd16,  9'd341},{  1'b0, 1'b0,  8'd14,   9'd82},{  1'b0, 1'b0,   8'd8,   9'd62},{  1'b0, 1'b0,   8'd2,  9'd242},{  1'b0, 1'b1,   8'd1,  9'd138},
{  1'b0, 1'b0, 8'd175,    9'd0},{  1'b0, 1'b0, 8'd174,    9'd0},{  1'b0, 1'b0, 8'd139,    9'd0},{  1'b0, 1'b0, 8'd110,  9'd342},{  1'b0, 1'b0, 8'd109,  9'd301},{  1'b0, 1'b0, 8'd103,    9'd0},{  1'b0, 1'b0,  8'd80,  9'd107},{  1'b0, 1'b0,  8'd72,  9'd156},{  1'b0, 1'b0,  8'd71,  9'd111},{  1'b0, 1'b0,  8'd67,    9'd0},{  1'b0, 1'b0,  8'd37,  9'd155},{  1'b0, 1'b0,  8'd34,  9'd354},{  1'b0, 1'b0,  8'd31,    9'd0},{  1'b0, 1'b0,  8'd23,  9'd340},{  1'b0, 1'b0,  8'd13,  9'd145},{  1'b0, 1'b0,   8'd8,  9'd219},{  1'b0, 1'b0,   8'd0,  9'd154},{  1'b0, 1'b1,   8'd0,  9'd348},
{  1'b0, 1'b0, 8'd176,    9'd0},{  1'b0, 1'b0, 8'd175,    9'd0},{  1'b0, 1'b0, 8'd141,   9'd74},{  1'b0, 1'b0, 8'd140,    9'd0},{  1'b0, 1'b0, 8'd132,  9'd240},{  1'b0, 1'b0, 8'd104,    9'd0},{  1'b0, 1'b0,  8'd91,   9'd70},{  1'b0, 1'b0,  8'd82,  9'd165},{  1'b0, 1'b0,  8'd68,    9'd0},{  1'b0, 1'b0,  8'd48,  9'd210},{  1'b0, 1'b0,  8'd43,  9'd142},{  1'b0, 1'b0,  8'd32,    9'd0},{  1'b0, 1'b0,  8'd31,  9'd252},{  1'b0, 1'b0,  8'd24,  9'd189},{  1'b0, 1'b0,  8'd14,  9'd264},{  1'b0, 1'b0,  8'd11,  9'd312},{  1'b0, 1'b0,   8'd8,  9'd195},{  1'b0, 1'b1,   8'd1,   9'd85},
{  1'b0, 1'b0, 8'd177,    9'd0},{  1'b0, 1'b0, 8'd176,    9'd0},{  1'b0, 1'b0, 8'd141,    9'd0},{  1'b0, 1'b0, 8'd140,   9'd68},{  1'b0, 1'b0, 8'd114,   9'd83},{  1'b0, 1'b0, 8'd105,    9'd0},{  1'b0, 1'b0, 8'd103,  9'd174},{  1'b0, 1'b0,  8'd95,   9'd58},{  1'b0, 1'b0,  8'd69,    9'd0},{  1'b0, 1'b0,  8'd66,  9'd327},{  1'b0, 1'b0,  8'd36,  9'd317},{  1'b0, 1'b0,  8'd33,    9'd0},{  1'b0, 1'b0,  8'd16,   9'd48},{  1'b0, 1'b0,  8'd12,  9'd286},{  1'b0, 1'b0,   8'd9,  9'd107},{  1'b0, 1'b0,   8'd4,   9'd14},{  1'b0, 1'b0,   8'd3,   9'd78},{  1'b0, 1'b1,   8'd2,   9'd59},
{  1'b0, 1'b0, 8'd178,    9'd0},{  1'b0, 1'b0, 8'd177,    9'd0},{  1'b0, 1'b0, 8'd142,    9'd0},{  1'b0, 1'b0, 8'd126,  9'd189},{  1'b0, 1'b0, 8'd115,   9'd57},{  1'b0, 1'b0, 8'd106,    9'd0},{  1'b0, 1'b0,  8'd84,  9'd102},{  1'b0, 1'b0,  8'd73,   9'd51},{  1'b0, 1'b0,  8'd70,    9'd0},{  1'b0, 1'b0,  8'd59,  9'd243},{  1'b0, 1'b0,  8'd37,  9'd207},{  1'b0, 1'b0,  8'd34,    9'd0},{  1'b0, 1'b0,  8'd32,  9'd203},{  1'b0, 1'b0,  8'd18,  9'd116},{  1'b0, 1'b0,  8'd10,  9'd220},{  1'b0, 1'b0,   8'd9,  9'd103},{  1'b0, 1'b0,   8'd4,  9'd117},{  1'b0, 1'b1,   8'd3,  9'd231},
{  1'b0, 1'b0, 8'd179,    9'd0},{  1'b0, 1'b0, 8'd178,    9'd0},{  1'b0, 1'b0, 8'd143,    9'd0},{  1'b0, 1'b0, 8'd135,  9'd336},{  1'b0, 1'b0, 8'd108,  9'd273},{  1'b0, 1'b0, 8'd107,    9'd0},{  1'b0, 1'b0, 8'd102,  9'd226},{  1'b0, 1'b0,  8'd91,   9'd56},{  1'b0, 1'b0,  8'd71,    9'd0},{  1'b0, 1'b0,  8'd71,   9'd31},{  1'b0, 1'b0,  8'd38,  9'd119},{  1'b0, 1'b0,  8'd35,    9'd0},{  1'b0, 1'b0,  8'd23,  9'd107},{  1'b0, 1'b0,  8'd12,   9'd57},{  1'b0, 1'b0,  8'd10,  9'd239},{  1'b0, 1'b0,   8'd4,  9'd312},{  1'b0, 1'b0,   8'd3,   9'd74},{  1'b0, 1'b1,   8'd1,  9'd213}
};
localparam bit [18 : 0] cLARGE_HS_V_TAB_4BY5_PACKED[cLARGE_HS_TAB_4BY5_PACKED_SIZE] = '{
{8'd179, 1'b0,   10'd0},{8'd179, 1'b1, 10'd630},
{8'd178, 1'b0, 10'd612},{8'd178, 1'b1, 10'd631},
{8'd177, 1'b0, 10'd594},{8'd177, 1'b1, 10'd613},
{8'd176, 1'b0, 10'd576},{8'd176, 1'b1, 10'd595},
{8'd175, 1'b0, 10'd558},{8'd175, 1'b1, 10'd577},
{8'd174, 1'b0, 10'd540},{8'd174, 1'b1, 10'd559},
{8'd173, 1'b0, 10'd522},{8'd173, 1'b1, 10'd541},
{8'd172, 1'b0, 10'd504},{8'd172, 1'b1, 10'd523},
{8'd171, 1'b0, 10'd486},{8'd171, 1'b1, 10'd505},
{8'd170, 1'b0, 10'd468},{8'd170, 1'b1, 10'd487},
{8'd169, 1'b0, 10'd450},{8'd169, 1'b1, 10'd469},
{8'd168, 1'b0, 10'd432},{8'd168, 1'b1, 10'd451},
{8'd167, 1'b0, 10'd414},{8'd167, 1'b1, 10'd433},
{8'd166, 1'b0, 10'd396},{8'd166, 1'b1, 10'd415},
{8'd165, 1'b0, 10'd378},{8'd165, 1'b1, 10'd397},
{8'd164, 1'b0, 10'd360},{8'd164, 1'b1, 10'd379},
{8'd163, 1'b0, 10'd342},{8'd163, 1'b1, 10'd361},
{8'd162, 1'b0, 10'd324},{8'd162, 1'b1, 10'd343},
{8'd161, 1'b0, 10'd306},{8'd161, 1'b1, 10'd325},
{8'd160, 1'b0, 10'd288},{8'd160, 1'b1, 10'd307},
{8'd159, 1'b0, 10'd270},{8'd159, 1'b1, 10'd289},
{8'd158, 1'b0, 10'd252},{8'd158, 1'b1, 10'd271},
{8'd157, 1'b0, 10'd234},{8'd157, 1'b1, 10'd253},
{8'd156, 1'b0, 10'd216},{8'd156, 1'b1, 10'd235},
{8'd155, 1'b0, 10'd198},{8'd155, 1'b1, 10'd217},
{8'd154, 1'b0, 10'd180},{8'd154, 1'b1, 10'd199},
{8'd153, 1'b0, 10'd162},{8'd153, 1'b1, 10'd181},
{8'd152, 1'b0, 10'd144},{8'd152, 1'b1, 10'd163},
{8'd151, 1'b0, 10'd126},{8'd151, 1'b1, 10'd145},
{8'd150, 1'b0, 10'd108},{8'd150, 1'b1, 10'd127},
{8'd149, 1'b0,  10'd90},{8'd149, 1'b1, 10'd109},
{8'd148, 1'b0,  10'd72},{8'd148, 1'b1,  10'd91},
{8'd147, 1'b0,  10'd54},{8'd147, 1'b1,  10'd73},
{8'd146, 1'b0,  10'd36},{8'd146, 1'b1,  10'd55},
{8'd145, 1'b0,  10'd18},{8'd145, 1'b1,  10'd37},
{8'd144, 1'b0,   10'd1},{8'd144, 1'b1,  10'd19},
{8'd143, 1'b0, 10'd164},{8'd143, 1'b0, 10'd290},{8'd143, 1'b1, 10'd632},
{8'd142, 1'b0, 10'd488},{8'd142, 1'b0, 10'd524},{8'd142, 1'b1, 10'd614},
{8'd141, 1'b0, 10'd291},{8'd141, 1'b0, 10'd578},{8'd141, 1'b1, 10'd596},
{8'd140, 1'b0, 10'd489},{8'd140, 1'b0, 10'd579},{8'd140, 1'b1, 10'd597},
{8'd139, 1'b0,   10'd2},{8'd139, 1'b0, 10'd362},{8'd139, 1'b1, 10'd560},
{8'd138, 1'b0, 10'd398},{8'd138, 1'b0, 10'd525},{8'd138, 1'b1, 10'd542},
{8'd137, 1'b0, 10'd416},{8'd137, 1'b0, 10'd434},{8'd137, 1'b1, 10'd526},
{8'd136, 1'b0, 10'd128},{8'd136, 1'b0, 10'd200},{8'd136, 1'b1, 10'd506},
{8'd135, 1'b0, 10'd110},{8'd135, 1'b0, 10'd490},{8'd135, 1'b1, 10'd633},
{8'd134, 1'b0,  10'd74},{8'd134, 1'b0, 10'd218},{8'd134, 1'b1, 10'd470},
{8'd133, 1'b0, 10'd146},{8'd133, 1'b0, 10'd452},{8'd133, 1'b1, 10'd453},
{8'd132, 1'b0, 10'd111},{8'd132, 1'b0, 10'd435},{8'd132, 1'b1, 10'd580},
{8'd131, 1'b0, 10'd236},{8'd131, 1'b0, 10'd380},{8'd131, 1'b1, 10'd417},
{8'd130, 1'b0, 10'd254},{8'd130, 1'b0, 10'd399},{8'd130, 1'b1, 10'd507},
{8'd129, 1'b0,  10'd56},{8'd129, 1'b0,  10'd92},{8'd129, 1'b1, 10'd381},
{8'd128, 1'b0,  10'd57},{8'd128, 1'b0,  10'd93},{8'd128, 1'b1, 10'd363},
{8'd127, 1'b0, 10'd255},{8'd127, 1'b0, 10'd326},{8'd127, 1'b1, 10'd344},
{8'd126, 1'b0, 10'd201},{8'd126, 1'b0, 10'd327},{8'd126, 1'b1, 10'd615},
{8'd125, 1'b0,   10'd3},{8'd125, 1'b0,  10'd38},{8'd125, 1'b1, 10'd308},
{8'd124, 1'b0, 10'd292},{8'd124, 1'b0, 10'd309},{8'd124, 1'b1, 10'd310},
{8'd123, 1'b0, 10'd165},{8'd123, 1'b0, 10'd272},{8'd123, 1'b1, 10'd328},
{8'd122, 1'b0,  10'd75},{8'd122, 1'b0, 10'd182},{8'd122, 1'b1, 10'd256},
{8'd121, 1'b0,  10'd20},{8'd121, 1'b0, 10'd237},{8'd121, 1'b1, 10'd273},
{8'd120, 1'b0, 10'd183},{8'd120, 1'b0, 10'd219},{8'd120, 1'b1, 10'd508},
{8'd119, 1'b0, 10'd202},{8'd119, 1'b0, 10'd345},{8'd119, 1'b1, 10'd471},
{8'd118, 1'b0,  10'd21},{8'd118, 1'b0,  10'd39},{8'd118, 1'b1, 10'd184},
{8'd117, 1'b0, 10'd166},{8'd117, 1'b0, 10'd364},{8'd117, 1'b1, 10'd454},
{8'd116, 1'b0, 10'd129},{8'd116, 1'b0, 10'd147},{8'd116, 1'b1, 10'd382},
{8'd115, 1'b0, 10'd130},{8'd115, 1'b0, 10'd472},{8'd115, 1'b1, 10'd616},
{8'd114, 1'b0, 10'd112},{8'd114, 1'b0, 10'd543},{8'd114, 1'b1, 10'd598},
{8'd113, 1'b0,  10'd94},{8'd113, 1'b0, 10'd220},{8'd113, 1'b1, 10'd418},
{8'd112, 1'b0,  10'd76},{8'd112, 1'b0, 10'd148},{8'd112, 1'b1, 10'd544},
{8'd111, 1'b0,  10'd58},{8'd111, 1'b0, 10'd274},{8'd111, 1'b1, 10'd400},
{8'd110, 1'b0,  10'd40},{8'd110, 1'b0, 10'd346},{8'd110, 1'b1, 10'd561},
{8'd109, 1'b0,  10'd22},{8'd109, 1'b0, 10'd436},{8'd109, 1'b1, 10'd562},
{8'd108, 1'b0,   10'd4},{8'd108, 1'b0, 10'd238},{8'd108, 1'b1, 10'd634},
{8'd107, 1'b0, 10'd275},{8'd107, 1'b0, 10'd365},{8'd107, 1'b1, 10'd635},
{8'd106, 1'b0,  10'd41},{8'd106, 1'b0, 10'd167},{8'd106, 1'b1, 10'd617},
{8'd105, 1'b0,  10'd95},{8'd105, 1'b0, 10'd545},{8'd105, 1'b1, 10'd599},
{8'd104, 1'b0,  10'd77},{8'd104, 1'b0, 10'd329},{8'd104, 1'b1, 10'd581},
{8'd103, 1'b0, 10'd437},{8'd103, 1'b0, 10'd563},{8'd103, 1'b1, 10'd600},
{8'd102, 1'b0, 10'd455},{8'd102, 1'b0, 10'd546},{8'd102, 1'b1, 10'd636},
{8'd101, 1'b0, 10'd419},{8'd101, 1'b0, 10'd509},{8'd101, 1'b1, 10'd527},
{8'd100, 1'b0, 10'd149},{8'd100, 1'b0, 10'd293},{8'd100, 1'b1, 10'd510},
{ 8'd99, 1'b0, 10'd168},{ 8'd99, 1'b0, 10'd276},{ 8'd99, 1'b1, 10'd491},
{ 8'd98, 1'b0,  10'd23},{ 8'd98, 1'b0, 10'd473},{ 8'd98, 1'b1, 10'd528},
{ 8'd97, 1'b0,  10'd96},{ 8'd97, 1'b0, 10'd347},{ 8'd97, 1'b1, 10'd456},
{ 8'd96, 1'b0,  10'd24},{ 8'd96, 1'b0, 10'd311},{ 8'd96, 1'b1, 10'd438},
{ 8'd95, 1'b0, 10'd420},{ 8'd95, 1'b0, 10'd457},{ 8'd95, 1'b1, 10'd601},
{ 8'd94, 1'b0,  10'd59},{ 8'd94, 1'b0, 10'd401},{ 8'd94, 1'b1, 10'd547},
{ 8'd93, 1'b0, 10'd330},{ 8'd93, 1'b0, 10'd383},{ 8'd93, 1'b1, 10'd511},
{ 8'd92, 1'b0, 10'd185},{ 8'd92, 1'b0, 10'd366},{ 8'd92, 1'b1, 10'd384},
{ 8'd91, 1'b0, 10'd348},{ 8'd91, 1'b0, 10'd582},{ 8'd91, 1'b1, 10'd637},
{ 8'd90, 1'b0, 10'd203},{ 8'd90, 1'b0, 10'd331},{ 8'd90, 1'b1, 10'd492},
{ 8'd89, 1'b0, 10'd312},{ 8'd89, 1'b0, 10'd421},{ 8'd89, 1'b1, 10'd529},
{ 8'd88, 1'b0, 10'd113},{ 8'd88, 1'b0, 10'd114},{ 8'd88, 1'b1, 10'd294},
{ 8'd87, 1'b0, 10'd257},{ 8'd87, 1'b0, 10'd277},{ 8'd87, 1'b1, 10'd474},
{ 8'd86, 1'b0,   10'd5},{ 8'd86, 1'b0, 10'd131},{ 8'd86, 1'b1, 10'd258},
{ 8'd85, 1'b0, 10'd221},{ 8'd85, 1'b0, 10'd239},{ 8'd85, 1'b1, 10'd493},
{ 8'd84, 1'b0,  10'd78},{ 8'd84, 1'b0, 10'd222},{ 8'd84, 1'b1, 10'd618},
{ 8'd83, 1'b0, 10'd204},{ 8'd83, 1'b0, 10'd240},{ 8'd83, 1'b1, 10'd259},
{ 8'd82, 1'b0, 10'd186},{ 8'd82, 1'b0, 10'd349},{ 8'd82, 1'b1, 10'd583},
{ 8'd81, 1'b0,   10'd6},{ 8'd81, 1'b0, 10'd169},{ 8'd81, 1'b1, 10'd187},
{ 8'd80, 1'b0, 10'd150},{ 8'd80, 1'b0, 10'd223},{ 8'd80, 1'b1, 10'd564},
{ 8'd79, 1'b0, 10'd132},{ 8'd79, 1'b0, 10'd313},{ 8'd79, 1'b1, 10'd367},
{ 8'd78, 1'b0,  10'd42},{ 8'd78, 1'b0, 10'd115},{ 8'd78, 1'b1, 10'd295},
{ 8'd77, 1'b0,  10'd97},{ 8'd77, 1'b0, 10'd151},{ 8'd77, 1'b1, 10'd385},
{ 8'd76, 1'b0,  10'd79},{ 8'd76, 1'b0, 10'd241},{ 8'd76, 1'b1, 10'd402},
{ 8'd75, 1'b0,  10'd60},{ 8'd75, 1'b0, 10'd205},{ 8'd75, 1'b1, 10'd403},
{ 8'd74, 1'b0,  10'd43},{ 8'd74, 1'b0, 10'd439},{ 8'd74, 1'b1, 10'd475},
{ 8'd73, 1'b0,  10'd25},{ 8'd73, 1'b0, 10'd133},{ 8'd73, 1'b1, 10'd619},
{ 8'd72, 1'b0,   10'd7},{ 8'd72, 1'b0,  10'd61},{ 8'd72, 1'b1, 10'd565},
{ 8'd71, 1'b0, 10'd566},{ 8'd71, 1'b0, 10'd638},{ 8'd71, 1'b1, 10'd639},
{ 8'd70, 1'b0, 10'd152},{ 8'd70, 1'b0, 10'd242},{ 8'd70, 1'b1, 10'd620},
{ 8'd69, 1'b0, 10'd260},{ 8'd69, 1'b0, 10'd296},{ 8'd69, 1'b1, 10'd602},
{ 8'd68, 1'b0, 10'd278},{ 8'd68, 1'b0, 10'd314},{ 8'd68, 1'b1, 10'd584},
{ 8'd67, 1'b0,  10'd44},{ 8'd67, 1'b0, 10'd243},{ 8'd67, 1'b1, 10'd567},
{ 8'd66, 1'b0, 10'd494},{ 8'd66, 1'b0, 10'd548},{ 8'd66, 1'b1, 10'd603},
{ 8'd65, 1'b0, 10'd188},{ 8'd65, 1'b0, 10'd206},{ 8'd65, 1'b1, 10'd530},
{ 8'd64, 1'b0, 10'd458},{ 8'd64, 1'b0, 10'd459},{ 8'd64, 1'b1, 10'd512},
{ 8'd63, 1'b0,  10'd26},{ 8'd63, 1'b0, 10'd134},{ 8'd63, 1'b1, 10'd495},
{ 8'd62, 1'b0, 10'd261},{ 8'd62, 1'b0, 10'd297},{ 8'd62, 1'b1, 10'd476},
{ 8'd61, 1'b0, 10'd224},{ 8'd61, 1'b0, 10'd422},{ 8'd61, 1'b1, 10'd460},
{ 8'd60, 1'b0, 10'd170},{ 8'd60, 1'b0, 10'd386},{ 8'd60, 1'b1, 10'd440},
{ 8'd59, 1'b0, 10'd332},{ 8'd59, 1'b0, 10'd423},{ 8'd59, 1'b1, 10'd621},
{ 8'd58, 1'b0,  10'd62},{ 8'd58, 1'b0, 10'd404},{ 8'd58, 1'b1, 10'd513},
{ 8'd57, 1'b0, 10'd116},{ 8'd57, 1'b0, 10'd279},{ 8'd57, 1'b1, 10'd387},
{ 8'd56, 1'b0, 10'd207},{ 8'd56, 1'b0, 10'd368},{ 8'd56, 1'b1, 10'd388},
{ 8'd55, 1'b0, 10'd350},{ 8'd55, 1'b0, 10'd441},{ 8'd55, 1'b1, 10'd531},
{ 8'd54, 1'b0,  10'd80},{ 8'd54, 1'b0, 10'd333},{ 8'd54, 1'b1, 10'd351},
{ 8'd53, 1'b0, 10'd315},{ 8'd53, 1'b0, 10'd334},{ 8'd53, 1'b1, 10'd532},
{ 8'd52, 1'b0, 10'd153},{ 8'd52, 1'b0, 10'd298},{ 8'd52, 1'b1, 10'd369},
{ 8'd51, 1'b0,  10'd98},{ 8'd51, 1'b0, 10'd280},{ 8'd51, 1'b1, 10'd549},
{ 8'd50, 1'b0, 10'd262},{ 8'd50, 1'b0, 10'd442},{ 8'd50, 1'b1, 10'd477},
{ 8'd49, 1'b0,   10'd8},{ 8'd49, 1'b0,  10'd81},{ 8'd49, 1'b1, 10'd244},
{ 8'd48, 1'b0,  10'd45},{ 8'd48, 1'b0, 10'd225},{ 8'd48, 1'b1, 10'd585},
{ 8'd47, 1'b0, 10'd189},{ 8'd47, 1'b0, 10'd208},{ 8'd47, 1'b1, 10'd550},
{ 8'd46, 1'b0, 10'd190},{ 8'd46, 1'b0, 10'd226},{ 8'd46, 1'b1, 10'd316},
{ 8'd45, 1'b0, 10'd135},{ 8'd45, 1'b0, 10'd171},{ 8'd45, 1'b1, 10'd405},
{ 8'd44, 1'b0,  10'd99},{ 8'd44, 1'b0, 10'd154},{ 8'd44, 1'b1, 10'd496},
{ 8'd43, 1'b0, 10'd136},{ 8'd43, 1'b0, 10'd406},{ 8'd43, 1'b1, 10'd586},
{ 8'd42, 1'b0, 10'd117},{ 8'd42, 1'b0, 10'd118},{ 8'd42, 1'b1, 10'd424},
{ 8'd41, 1'b0,  10'd27},{ 8'd41, 1'b0, 10'd100},{ 8'd41, 1'b1, 10'd514},
{ 8'd40, 1'b0,  10'd63},{ 8'd40, 1'b0,  10'd82},{ 8'd40, 1'b1, 10'd478},
{ 8'd39, 1'b0,   10'd9},{ 8'd39, 1'b0,  10'd64},{ 8'd39, 1'b1, 10'd370},
{ 8'd38, 1'b0,  10'd46},{ 8'd38, 1'b0, 10'd352},{ 8'd38, 1'b1, 10'd640},
{ 8'd37, 1'b0,  10'd28},{ 8'd37, 1'b0, 10'd568},{ 8'd37, 1'b1, 10'd622},
{ 8'd36, 1'b0,  10'd10},{ 8'd36, 1'b0, 10'd172},{ 8'd36, 1'b1, 10'd604},
{ 8'd35, 1'b0, 10'd335},{ 8'd35, 1'b0, 10'd551},{ 8'd35, 1'b1, 10'd641},
{ 8'd34, 1'b0, 10'd425},{ 8'd34, 1'b0, 10'd569},{ 8'd34, 1'b1, 10'd623},
{ 8'd33, 1'b0,  10'd29},{ 8'd33, 1'b0, 10'd209},{ 8'd33, 1'b1, 10'd605},
{ 8'd32, 1'b0, 10'd263},{ 8'd32, 1'b0, 10'd587},{ 8'd32, 1'b1, 10'd624},
{ 8'd31, 1'b0,  10'd83},{ 8'd31, 1'b0, 10'd570},{ 8'd31, 1'b1, 10'd588},
{ 8'd30, 1'b0,  10'd84},{ 8'd30, 1'b0, 10'd227},{ 8'd30, 1'b1, 10'd552},
{ 8'd29, 1'b0, 10'd245},{ 8'd29, 1'b0, 10'd371},{ 8'd29, 1'b1, 10'd533},
{ 8'd28, 1'b0, 10'd461},{ 8'd28, 1'b0, 10'd515},{ 8'd28, 1'b1, 10'd534},
{ 8'd27, 1'b0,  10'd30},{ 8'd27, 1'b0, 10'd119},{ 8'd27, 1'b1, 10'd497},
{ 8'd26, 1'b0, 10'd173},{ 8'd26, 1'b0, 10'd389},{ 8'd26, 1'b1, 10'd479},
{ 8'd25, 1'b0,  10'd11},{ 8'd25, 1'b0, 10'd191},{ 8'd25, 1'b1, 10'd462},
{ 8'd24, 1'b0, 10'd443},{ 8'd24, 1'b0, 10'd516},{ 8'd24, 1'b1, 10'd589},
{ 8'd23, 1'b0, 10'd426},{ 8'd23, 1'b0, 10'd571},{ 8'd23, 1'b1, 10'd642},
{ 8'd22, 1'b0, 10'd101},{ 8'd22, 1'b0, 10'd264},{ 8'd22, 1'b1, 10'd407},
{ 8'd21, 1'b0,  10'd47},{ 8'd21, 1'b0, 10'd353},{ 8'd21, 1'b1, 10'd390},
{ 8'd20, 1'b0, 10'd155},{ 8'd20, 1'b0, 10'd372},{ 8'd20, 1'b1, 10'd480},
{ 8'd19, 1'b0,  10'd48},{ 8'd19, 1'b0, 10'd137},{ 8'd19, 1'b1, 10'd354},
{ 8'd18, 1'b0,  10'd65},{ 8'd18, 1'b0, 10'd336},{ 8'd18, 1'b1, 10'd625},
{ 8'd17, 1'b0,  10'd12},{ 8'd17, 1'b0,  10'd31},{ 8'd17, 1'b0, 10'd265},{ 8'd17, 1'b0, 10'd299},{ 8'd17, 1'b0, 10'd317},{ 8'd17, 1'b0, 10'd318},{ 8'd17, 1'b0, 10'd373},{ 8'd17, 1'b0, 10'd391},{ 8'd17, 1'b0, 10'd463},{ 8'd17, 1'b0, 10'd464},{ 8'd17, 1'b1, 10'd517},
{ 8'd16, 1'b0, 10'd102},{ 8'd16, 1'b0, 10'd246},{ 8'd16, 1'b0, 10'd300},{ 8'd16, 1'b0, 10'd337},{ 8'd16, 1'b0, 10'd355},{ 8'd16, 1'b0, 10'd408},{ 8'd16, 1'b0, 10'd409},{ 8'd16, 1'b0, 10'd410},{ 8'd16, 1'b0, 10'd535},{ 8'd16, 1'b0, 10'd553},{ 8'd16, 1'b1, 10'd606},
{ 8'd15, 1'b0,  10'd13},{ 8'd15, 1'b0,  10'd14},{ 8'd15, 1'b0,  10'd66},{ 8'd15, 1'b0,  10'd85},{ 8'd15, 1'b0, 10'd210},{ 8'd15, 1'b0, 10'd211},{ 8'd15, 1'b0, 10'd266},{ 8'd15, 1'b0, 10'd281},{ 8'd15, 1'b0, 10'd301},{ 8'd15, 1'b0, 10'd444},{ 8'd15, 1'b1, 10'd498},
{ 8'd14, 1'b0,  10'd32},{ 8'd14, 1'b0, 10'd138},{ 8'd14, 1'b0, 10'd156},{ 8'd14, 1'b0, 10'd267},{ 8'd14, 1'b0, 10'd374},{ 8'd14, 1'b0, 10'd392},{ 8'd14, 1'b0, 10'd393},{ 8'd14, 1'b0, 10'd465},{ 8'd14, 1'b0, 10'd536},{ 8'd14, 1'b0, 10'd554},{ 8'd14, 1'b1, 10'd590},
{ 8'd13, 1'b0, 10'd103},{ 8'd13, 1'b0, 10'd120},{ 8'd13, 1'b0, 10'd174},{ 8'd13, 1'b0, 10'd192},{ 8'd13, 1'b0, 10'd247},{ 8'd13, 1'b0, 10'd394},{ 8'd13, 1'b0, 10'd466},{ 8'd13, 1'b0, 10'd481},{ 8'd13, 1'b0, 10'd499},{ 8'd13, 1'b0, 10'd537},{ 8'd13, 1'b1, 10'd572},
{ 8'd12, 1'b0,  10'd15},{ 8'd12, 1'b0,  10'd49},{ 8'd12, 1'b0, 10'd193},{ 8'd12, 1'b0, 10'd194},{ 8'd12, 1'b0, 10'd212},{ 8'd12, 1'b0, 10'd228},{ 8'd12, 1'b0, 10'd282},{ 8'd12, 1'b0, 10'd338},{ 8'd12, 1'b0, 10'd538},{ 8'd12, 1'b0, 10'd607},{ 8'd12, 1'b1, 10'd643},
{ 8'd11, 1'b0,  10'd67},{ 8'd11, 1'b0, 10'd121},{ 8'd11, 1'b0, 10'd122},{ 8'd11, 1'b0, 10'd213},{ 8'd11, 1'b0, 10'd229},{ 8'd11, 1'b0, 10'd268},{ 8'd11, 1'b0, 10'd283},{ 8'd11, 1'b0, 10'd302},{ 8'd11, 1'b0, 10'd356},{ 8'd11, 1'b0, 10'd445},{ 8'd11, 1'b1, 10'd591},
{ 8'd10, 1'b0,  10'd33},{ 8'd10, 1'b0,  10'd50},{ 8'd10, 1'b0, 10'd139},{ 8'd10, 1'b0, 10'd140},{ 8'd10, 1'b0, 10'd157},{ 8'd10, 1'b0, 10'd195},{ 8'd10, 1'b0, 10'd230},{ 8'd10, 1'b0, 10'd482},{ 8'd10, 1'b0, 10'd500},{ 8'd10, 1'b0, 10'd626},{ 8'd10, 1'b1, 10'd644},
{  8'd9, 1'b0,  10'd34},{  8'd9, 1'b0,  10'd68},{  8'd9, 1'b0, 10'd104},{  8'd9, 1'b0, 10'd158},{  8'd9, 1'b0, 10'd175},{  8'd9, 1'b0, 10'd248},{  8'd9, 1'b0, 10'd339},{  8'd9, 1'b0, 10'd483},{  8'd9, 1'b0, 10'd501},{  8'd9, 1'b0, 10'd608},{  8'd9, 1'b1, 10'd627},
{  8'd8, 1'b0, 10'd123},{  8'd8, 1'b0, 10'd159},{  8'd8, 1'b0, 10'd160},{  8'd8, 1'b0, 10'd214},{  8'd8, 1'b0, 10'd215},{  8'd8, 1'b0, 10'd319},{  8'd8, 1'b0, 10'd340},{  8'd8, 1'b0, 10'd502},{  8'd8, 1'b0, 10'd555},{  8'd8, 1'b0, 10'd573},{  8'd8, 1'b1, 10'd592},
{  8'd7, 1'b0,  10'd51},{  8'd7, 1'b0,  10'd86},{  8'd7, 1'b0, 10'd124},{  8'd7, 1'b0, 10'd141},{  8'd7, 1'b0, 10'd249},{  8'd7, 1'b0, 10'd269},{  8'd7, 1'b0, 10'd284},{  8'd7, 1'b0, 10'd285},{  8'd7, 1'b0, 10'd427},{  8'd7, 1'b0, 10'd428},{  8'd7, 1'b1, 10'd429},
{  8'd6, 1'b0,  10'd16},{  8'd6, 1'b0,  10'd87},{  8'd6, 1'b0, 10'd125},{  8'd6, 1'b0, 10'd142},{  8'd6, 1'b0, 10'd303},{  8'd6, 1'b0, 10'd320},{  8'd6, 1'b0, 10'd411},{  8'd6, 1'b0, 10'd412},{  8'd6, 1'b0, 10'd484},{  8'd6, 1'b0, 10'd503},{  8'd6, 1'b1, 10'd518},
{  8'd5, 1'b0,  10'd52},{  8'd5, 1'b0,  10'd69},{  8'd5, 1'b0,  10'd70},{  8'd5, 1'b0, 10'd105},{  8'd5, 1'b0, 10'd106},{  8'd5, 1'b0, 10'd286},{  8'd5, 1'b0, 10'd304},{  8'd5, 1'b0, 10'd357},{  8'd5, 1'b0, 10'd446},{  8'd5, 1'b0, 10'd447},{  8'd5, 1'b1, 10'd519},
{  8'd4, 1'b0,  10'd88},{  8'd4, 1'b0,  10'd89},{  8'd4, 1'b0, 10'd143},{  8'd4, 1'b0, 10'd196},{  8'd4, 1'b0, 10'd250},{  8'd4, 1'b0, 10'd358},{  8'd4, 1'b0, 10'd430},{  8'd4, 1'b0, 10'd431},{  8'd4, 1'b0, 10'd609},{  8'd4, 1'b0, 10'd628},{  8'd4, 1'b1, 10'd645},
{  8'd3, 1'b0,  10'd71},{  8'd3, 1'b0, 10'd197},{  8'd3, 1'b0, 10'd251},{  8'd3, 1'b0, 10'd287},{  8'd3, 1'b0, 10'd375},{  8'd3, 1'b0, 10'd467},{  8'd3, 1'b0, 10'd520},{  8'd3, 1'b0, 10'd521},{  8'd3, 1'b0, 10'd610},{  8'd3, 1'b0, 10'd629},{  8'd3, 1'b1, 10'd646},
{  8'd2, 1'b0,  10'd53},{  8'd2, 1'b0, 10'd176},{  8'd2, 1'b0, 10'd177},{  8'd2, 1'b0, 10'd231},{  8'd2, 1'b0, 10'd359},{  8'd2, 1'b0, 10'd376},{  8'd2, 1'b0, 10'd377},{  8'd2, 1'b0, 10'd448},{  8'd2, 1'b0, 10'd539},{  8'd2, 1'b0, 10'd556},{  8'd2, 1'b1, 10'd611},
{  8'd1, 1'b0,  10'd35},{  8'd1, 1'b0, 10'd178},{  8'd1, 1'b0, 10'd321},{  8'd1, 1'b0, 10'd322},{  8'd1, 1'b0, 10'd323},{  8'd1, 1'b0, 10'd395},{  8'd1, 1'b0, 10'd413},{  8'd1, 1'b0, 10'd485},{  8'd1, 1'b0, 10'd557},{  8'd1, 1'b0, 10'd593},{  8'd1, 1'b1, 10'd647},
{  8'd0, 1'b0,  10'd17},{  8'd0, 1'b0, 10'd107},{  8'd0, 1'b0, 10'd161},{  8'd0, 1'b0, 10'd179},{  8'd0, 1'b0, 10'd232},{  8'd0, 1'b0, 10'd233},{  8'd0, 1'b0, 10'd305},{  8'd0, 1'b0, 10'd341},{  8'd0, 1'b0, 10'd449},{  8'd0, 1'b0, 10'd574},{  8'd0, 1'b1, 10'd575}
};
localparam int          cLARGE_HS_TAB_5BY6_PACKED_SIZE = 660;
localparam bit [18 : 0] cLARGE_HS_TAB_5BY6_PACKED[cLARGE_HS_TAB_5BY6_PACKED_SIZE] = '{
{  1'b1, 1'b0, 8'd179,    9'd1},{  1'b0, 1'b0, 8'd150,    9'd0},{  1'b0, 1'b0, 8'd140,  9'd151},{  1'b0, 1'b0, 8'd136,  9'd111},{  1'b0, 1'b0, 8'd120,    9'd0},{  1'b0, 1'b0, 8'd118,  9'd161},{  1'b0, 1'b0,  8'd97,  9'd108},{  1'b0, 1'b0,  8'd90,    9'd0},{  1'b0, 1'b0,  8'd78,   9'd21},{  1'b0, 1'b0,  8'd72,  9'd280},{  1'b0, 1'b0,  8'd60,    9'd0},{  1'b0, 1'b0,  8'd54,  9'd280},{  1'b0, 1'b0,  8'd40,   9'd88},{  1'b0, 1'b0,  8'd30,    9'd0},{  1'b0, 1'b0,  8'd14,  9'd120},{  1'b0, 1'b0,  8'd14,   9'd19},{  1'b0, 1'b0,  8'd13,  9'd142},{  1'b0, 1'b0,   8'd9,  9'd128},{  1'b0, 1'b0,   8'd8,   9'd86},{  1'b0, 1'b0,   8'd6,  9'd332},{  1'b0, 1'b0,   8'd3,  9'd312},{  1'b0, 1'b1,   8'd0,    9'd0},
{  1'b0, 1'b0, 8'd151,    9'd0},{  1'b0, 1'b0, 8'd150,    9'd0},{  1'b0, 1'b0, 8'd148,   9'd71},{  1'b0, 1'b0, 8'd131,   9'd43},{  1'b0, 1'b0, 8'd121,    9'd0},{  1'b0, 1'b0, 8'd101,  9'd204},{  1'b0, 1'b0, 8'd100,  9'd191},{  1'b0, 1'b0,  8'd91,    9'd0},{  1'b0, 1'b0,  8'd69,  9'd211},{  1'b0, 1'b0,  8'd67,  9'd171},{  1'b0, 1'b0,  8'd61,    9'd0},{  1'b0, 1'b0,  8'd46,  9'd273},{  1'b0, 1'b0,  8'd31,    9'd0},{  1'b0, 1'b0,  8'd31,   9'd88},{  1'b0, 1'b0,  8'd19,  9'd284},{  1'b0, 1'b0,  8'd15,  9'd254},{  1'b0, 1'b0,  8'd13,  9'd223},{  1'b0, 1'b0,   8'd7,  9'd263},{  1'b0, 1'b0,   8'd2,  9'd103},{  1'b0, 1'b0,   8'd2,  9'd189},{  1'b0, 1'b0,   8'd1,    9'd0},{  1'b0, 1'b1,   8'd1,  9'd201},
{  1'b0, 1'b0, 8'd152,    9'd0},{  1'b0, 1'b0, 8'd151,    9'd0},{  1'b0, 1'b0, 8'd132,  9'd353},{  1'b0, 1'b0, 8'd130,  9'd204},{  1'b0, 1'b0, 8'd122,    9'd0},{  1'b0, 1'b0, 8'd116,   9'd12},{  1'b0, 1'b0,  8'd92,    9'd0},{  1'b0, 1'b0,  8'd91,  9'd120},{  1'b0, 1'b0,  8'd70,  9'd222},{  1'b0, 1'b0,  8'd65,  9'd155},{  1'b0, 1'b0,  8'd62,    9'd0},{  1'b0, 1'b0,  8'd56,  9'd168},{  1'b0, 1'b0,  8'd42,  9'd186},{  1'b0, 1'b0,  8'd32,    9'd0},{  1'b0, 1'b0,  8'd28,  9'd118},{  1'b0, 1'b0,  8'd27,  9'd169},{  1'b0, 1'b0,  8'd12,  9'd318},{  1'b0, 1'b0,  8'd12,  9'd245},{  1'b0, 1'b0,   8'd9,  9'd219},{  1'b0, 1'b0,   8'd5,  9'd135},{  1'b0, 1'b0,   8'd2,    9'd0},{  1'b0, 1'b1,   8'd0,   9'd97},
{  1'b0, 1'b0, 8'd153,    9'd0},{  1'b0, 1'b0, 8'd152,    9'd0},{  1'b0, 1'b0, 8'd148,  9'd156},{  1'b0, 1'b0, 8'd137,  9'd352},{  1'b0, 1'b0, 8'd123,    9'd0},{  1'b0, 1'b0, 8'd111,   9'd25},{  1'b0, 1'b0,  8'd93,    9'd0},{  1'b0, 1'b0,  8'd90,  9'd105},{  1'b0, 1'b0,  8'd79,   9'd12},{  1'b0, 1'b0,  8'd64,  9'd217},{  1'b0, 1'b0,  8'd63,    9'd0},{  1'b0, 1'b0,  8'd58,  9'd240},{  1'b0, 1'b0,  8'd34,  9'd250},{  1'b0, 1'b0,  8'd33,    9'd0},{  1'b0, 1'b0,  8'd17,  9'd243},{  1'b0, 1'b0,  8'd12,  9'd354},{  1'b0, 1'b0,  8'd11,  9'd353},{  1'b0, 1'b0,   8'd8,   9'd96},{  1'b0, 1'b0,   8'd5,  9'd123},{  1'b0, 1'b0,   8'd4,  9'd328},{  1'b0, 1'b0,   8'd3,    9'd0},{  1'b0, 1'b1,   8'd0,  9'd224},
{  1'b0, 1'b0, 8'd154,    9'd0},{  1'b0, 1'b0, 8'd153,    9'd0},{  1'b0, 1'b0, 8'd146,  9'd214},{  1'b0, 1'b0, 8'd137,  9'd142},{  1'b0, 1'b0, 8'd124,    9'd0},{  1'b0, 1'b0, 8'd113,   9'd87},{  1'b0, 1'b0, 8'd109,  9'd302},{  1'b0, 1'b0,  8'd94,    9'd0},{  1'b0, 1'b0,  8'd87,  9'd202},{  1'b0, 1'b0,  8'd77,   9'd95},{  1'b0, 1'b0,  8'd64,    9'd0},{  1'b0, 1'b0,  8'd55,   9'd13},{  1'b0, 1'b0,  8'd39,  9'd132},{  1'b0, 1'b0,  8'd34,    9'd0},{  1'b0, 1'b0,  8'd15,  9'd210},{  1'b0, 1'b0,  8'd11,   9'd13},{  1'b0, 1'b0,   8'd9,   9'd69},{  1'b0, 1'b0,   8'd9,  9'd103},{  1'b0, 1'b0,   8'd8,   9'd34},{  1'b0, 1'b0,   8'd5,  9'd238},{  1'b0, 1'b0,   8'd4,    9'd0},{  1'b0, 1'b1,   8'd4,  9'd261},
{  1'b0, 1'b0, 8'd155,    9'd0},{  1'b0, 1'b0, 8'd154,    9'd0},{  1'b0, 1'b0, 8'd147,  9'd125},{  1'b0, 1'b0, 8'd132,  9'd298},{  1'b0, 1'b0, 8'd125,    9'd0},{  1'b0, 1'b0, 8'd115,   9'd69},{  1'b0, 1'b0,  8'd95,    9'd0},{  1'b0, 1'b0,  8'd91,  9'd135},{  1'b0, 1'b0,  8'd89,   9'd96},{  1'b0, 1'b0,  8'd65,    9'd0},{  1'b0, 1'b0,  8'd63,  9'd353},{  1'b0, 1'b0,  8'd55,  9'd275},{  1'b0, 1'b0,  8'd48,  9'd110},{  1'b0, 1'b0,  8'd35,    9'd0},{  1'b0, 1'b0,  8'd13,  9'd125},{  1'b0, 1'b0,  8'd12,   9'd24},{  1'b0, 1'b0,   8'd8,   9'd73},{  1'b0, 1'b0,   8'd7,  9'd158},{  1'b0, 1'b0,   8'd5,    9'd0},{  1'b0, 1'b0,   8'd4,  9'd161},{  1'b0, 1'b0,   8'd2,  9'd339},{  1'b0, 1'b1,   8'd2,  9'd166},
{  1'b0, 1'b0, 8'd156,    9'd0},{  1'b0, 1'b0, 8'd155,    9'd0},{  1'b0, 1'b0, 8'd143,   9'd70},{  1'b0, 1'b0, 8'd129,  9'd322},{  1'b0, 1'b0, 8'd126,    9'd0},{  1'b0, 1'b0, 8'd111,  9'd244},{  1'b0, 1'b0, 8'd107,  9'd267},{  1'b0, 1'b0,  8'd96,    9'd0},{  1'b0, 1'b0,  8'd86,  9'd151},{  1'b0, 1'b0,  8'd73,  9'd305},{  1'b0, 1'b0,  8'd66,    9'd0},{  1'b0, 1'b0,  8'd45,  9'd150},{  1'b0, 1'b0,  8'd37,  9'd309},{  1'b0, 1'b0,  8'd36,    9'd0},{  1'b0, 1'b0,  8'd17,  9'd226},{  1'b0, 1'b0,  8'd11,  9'd121},{  1'b0, 1'b0,   8'd9,  9'd126},{  1'b0, 1'b0,   8'd7,  9'd139},{  1'b0, 1'b0,   8'd6,    9'd0},{  1'b0, 1'b0,   8'd6,  9'd277},{  1'b0, 1'b0,   8'd3,  9'd333},{  1'b0, 1'b1,   8'd0,  9'd107},
{  1'b0, 1'b0, 8'd157,    9'd0},{  1'b0, 1'b0, 8'd156,    9'd0},{  1'b0, 1'b0, 8'd127,    9'd0},{  1'b0, 1'b0, 8'd123,  9'd122},{  1'b0, 1'b0, 8'd120,  9'd261},{  1'b0, 1'b0, 8'd116,  9'd156},{  1'b0, 1'b0,  8'd97,    9'd0},{  1'b0, 1'b0,  8'd92,   9'd57},{  1'b0, 1'b0,  8'd83,  9'd192},{  1'b0, 1'b0,  8'd67,    9'd0},{  1'b0, 1'b0,  8'd62,    9'd2},{  1'b0, 1'b0,  8'd52,   9'd37},{  1'b0, 1'b0,  8'd47,  9'd205},{  1'b0, 1'b0,  8'd37,    9'd0},{  1'b0, 1'b0,  8'd27,   9'd35},{  1'b0, 1'b0,  8'd22,  9'd317},{  1'b0, 1'b0,   8'd7,    9'd0},{  1'b0, 1'b0,   8'd7,   9'd57},{  1'b0, 1'b0,   8'd7,   9'd52},{  1'b0, 1'b0,   8'd3,  9'd143},{  1'b0, 1'b0,   8'd2,  9'd242},{  1'b0, 1'b1,   8'd1,  9'd213},
{  1'b0, 1'b0, 8'd158,    9'd0},{  1'b0, 1'b0, 8'd157,    9'd0},{  1'b0, 1'b0, 8'd141,  9'd227},{  1'b0, 1'b0, 8'd130,  9'd236},{  1'b0, 1'b0, 8'd128,    9'd0},{  1'b0, 1'b0, 8'd100,  9'd262},{  1'b0, 1'b0,  8'd98,    9'd0},{  1'b0, 1'b0,  8'd94,  9'd263},{  1'b0, 1'b0,  8'd71,  9'd341},{  1'b0, 1'b0,  8'd68,    9'd0},{  1'b0, 1'b0,  8'd62,  9'd241},{  1'b0, 1'b0,  8'd56,  9'd211},{  1'b0, 1'b0,  8'd39,   9'd11},{  1'b0, 1'b0,  8'd38,    9'd0},{  1'b0, 1'b0,  8'd28,  9'd264},{  1'b0, 1'b0,  8'd22,  9'd342},{  1'b0, 1'b0,  8'd13,  9'd293},{  1'b0, 1'b0,  8'd12,  9'd252},{  1'b0, 1'b0,   8'd8,    9'd0},{  1'b0, 1'b0,   8'd3,  9'd335},{  1'b0, 1'b0,   8'd3,  9'd171},{  1'b0, 1'b1,   8'd1,  9'd299},
{  1'b0, 1'b0, 8'd159,    9'd0},{  1'b0, 1'b0, 8'd158,    9'd0},{  1'b0, 1'b0, 8'd133,  9'd120},{  1'b0, 1'b0, 8'd129,    9'd0},{  1'b0, 1'b0, 8'd121,   9'd56},{  1'b0, 1'b0, 8'd105,  9'd100},{  1'b0, 1'b0,  8'd99,    9'd0},{  1'b0, 1'b0,  8'd98,  9'd316},{  1'b0, 1'b0,  8'd82,  9'd302},{  1'b0, 1'b0,  8'd77,  9'd282},{  1'b0, 1'b0,  8'd69,    9'd0},{  1'b0, 1'b0,  8'd58,   9'd66},{  1'b0, 1'b0,  8'd53,  9'd187},{  1'b0, 1'b0,  8'd39,    9'd0},{  1'b0, 1'b0,  8'd13,  9'd247},{  1'b0, 1'b0,   8'd9,    9'd0},{  1'b0, 1'b0,   8'd8,   9'd56},{  1'b0, 1'b0,   8'd8,  9'd148},{  1'b0, 1'b0,   8'd6,  9'd173},{  1'b0, 1'b0,   8'd6,   9'd23},{  1'b0, 1'b0,   8'd4,   9'd79},{  1'b0, 1'b1,   8'd2,  9'd300},
{  1'b0, 1'b0, 8'd160,    9'd0},{  1'b0, 1'b0, 8'd159,    9'd0},{  1'b0, 1'b0, 8'd133,  9'd237},{  1'b0, 1'b0, 8'd130,    9'd0},{  1'b0, 1'b0, 8'd128,  9'd110},{  1'b0, 1'b0, 8'd117,  9'd331},{  1'b0, 1'b0, 8'd103,   9'd19},{  1'b0, 1'b0, 8'd100,    9'd0},{  1'b0, 1'b0,  8'd83,  9'd135},{  1'b0, 1'b0,  8'd76,   9'd56},{  1'b0, 1'b0,  8'd70,    9'd0},{  1'b0, 1'b0,  8'd49,   9'd51},{  1'b0, 1'b0,  8'd40,    9'd0},{  1'b0, 1'b0,  8'd34,  9'd313},{  1'b0, 1'b0,  8'd24,  9'd185},{  1'b0, 1'b0,  8'd18,  9'd198},{  1'b0, 1'b0,  8'd14,  9'd217},{  1'b0, 1'b0,  8'd10,    9'd0},{  1'b0, 1'b0,   8'd9,   9'd48},{  1'b0, 1'b0,   8'd4,  9'd102},{  1'b0, 1'b0,   8'd3,  9'd112},{  1'b0, 1'b1,   8'd0,   9'd85},
{  1'b0, 1'b0, 8'd161,    9'd0},{  1'b0, 1'b0, 8'd160,    9'd0},{  1'b0, 1'b0, 8'd145,   9'd72},{  1'b0, 1'b0, 8'd144,  9'd229},{  1'b0, 1'b0, 8'd131,    9'd0},{  1'b0, 1'b0, 8'd115,   9'd20},{  1'b0, 1'b0, 8'd101,    9'd0},{  1'b0, 1'b0,  8'd90,  9'd356},{  1'b0, 1'b0,  8'd89,   9'd68},{  1'b0, 1'b0,  8'd71,    9'd0},{  1'b0, 1'b0,  8'd63,  9'd294},{  1'b0, 1'b0,  8'd59,   9'd59},{  1'b0, 1'b0,  8'd45,  9'd116},{  1'b0, 1'b0,  8'd41,    9'd0},{  1'b0, 1'b0,  8'd13,  9'd238},{  1'b0, 1'b0,  8'd12,   9'd84},{  1'b0, 1'b0,  8'd11,    9'd0},{  1'b0, 1'b0,  8'd11,  9'd285},{  1'b0, 1'b0,   8'd6,  9'd344},{  1'b0, 1'b0,   8'd6,   9'd66},{  1'b0, 1'b0,   8'd5,  9'd262},{  1'b0, 1'b1,   8'd1,  9'd100},
{  1'b0, 1'b0, 8'd162,    9'd0},{  1'b0, 1'b0, 8'd161,    9'd0},{  1'b0, 1'b0, 8'd146,  9'd135},{  1'b0, 1'b0, 8'd135,  9'd268},{  1'b0, 1'b0, 8'd132,    9'd0},{  1'b0, 1'b0, 8'd102,    9'd0},{  1'b0, 1'b0, 8'd102,  9'd304},{  1'b0, 1'b0,  8'd98,  9'd222},{  1'b0, 1'b0,  8'd86,  9'd296},{  1'b0, 1'b0,  8'd81,  9'd223},{  1'b0, 1'b0,  8'd72,    9'd0},{  1'b0, 1'b0,  8'd46,  9'd139},{  1'b0, 1'b0,  8'd42,    9'd0},{  1'b0, 1'b0,  8'd37,   9'd56},{  1'b0, 1'b0,  8'd29,  9'd125},{  1'b0, 1'b0,  8'd12,    9'd0},{  1'b0, 1'b0,  8'd11,  9'd129},{  1'b0, 1'b0,  8'd10,  9'd315},{  1'b0, 1'b0,   8'd9,   9'd50},{  1'b0, 1'b0,   8'd7,  9'd358},{  1'b0, 1'b0,   8'd2,  9'd136},{  1'b0, 1'b1,   8'd0,  9'd145},
{  1'b0, 1'b0, 8'd163,    9'd0},{  1'b0, 1'b0, 8'd162,    9'd0},{  1'b0, 1'b0, 8'd144,  9'd129},{  1'b0, 1'b0, 8'd142,  9'd113},{  1'b0, 1'b0, 8'd133,    9'd0},{  1'b0, 1'b0, 8'd119,   9'd45},{  1'b0, 1'b0, 8'd103,    9'd0},{  1'b0, 1'b0, 8'd102,  9'd161},{  1'b0, 1'b0,  8'd88,  9'd196},{  1'b0, 1'b0,  8'd87,   9'd28},{  1'b0, 1'b0,  8'd73,    9'd0},{  1'b0, 1'b0,  8'd43,    9'd0},{  1'b0, 1'b0,  8'd43,  9'd317},{  1'b0, 1'b0,  8'd42,  9'd189},{  1'b0, 1'b0,  8'd13,    9'd0},{  1'b0, 1'b0,  8'd13,  9'd275},{  1'b0, 1'b0,  8'd12,   9'd54},{  1'b0, 1'b0,   8'd9,  9'd286},{  1'b0, 1'b0,   8'd7,  9'd229},{  1'b0, 1'b0,   8'd4,  9'd278},{  1'b0, 1'b0,   8'd1,  9'd310},{  1'b0, 1'b1,   8'd0,  9'd286},
{  1'b0, 1'b0, 8'd164,    9'd0},{  1'b0, 1'b0, 8'd163,    9'd0},{  1'b0, 1'b0, 8'd134,    9'd0},{  1'b0, 1'b0, 8'd127,  9'd131},{  1'b0, 1'b0, 8'd125,  9'd141},{  1'b0, 1'b0, 8'd117,  9'd289},{  1'b0, 1'b0, 8'd113,  9'd261},{  1'b0, 1'b0, 8'd104,    9'd0},{  1'b0, 1'b0,  8'd74,    9'd0},{  1'b0, 1'b0,  8'd71,  9'd320},{  1'b0, 1'b0,  8'd61,  9'd140},{  1'b0, 1'b0,  8'd59,  9'd172},{  1'b0, 1'b0,  8'd44,    9'd0},{  1'b0, 1'b0,  8'd32,   9'd92},{  1'b0, 1'b0,  8'd14,    9'd0},{  1'b0, 1'b0,  8'd12,    9'd2},{  1'b0, 1'b0,  8'd11,  9'd273},{  1'b0, 1'b0,   8'd9,  9'd181},{  1'b0, 1'b0,   8'd7,  9'd325},{  1'b0, 1'b0,   8'd6,   9'd43},{  1'b0, 1'b0,   8'd5,   9'd69},{  1'b0, 1'b1,   8'd3,   9'd14},
{  1'b0, 1'b0, 8'd165,    9'd0},{  1'b0, 1'b0, 8'd164,    9'd0},{  1'b0, 1'b0, 8'd136,   9'd96},{  1'b0, 1'b0, 8'd135,    9'd0},{  1'b0, 1'b0, 8'd126,  9'd341},{  1'b0, 1'b0, 8'd108,  9'd306},{  1'b0, 1'b0, 8'd106,    9'd6},{  1'b0, 1'b0, 8'd105,    9'd0},{  1'b0, 1'b0,  8'd80,  9'd137},{  1'b0, 1'b0,  8'd75,    9'd0},{  1'b0, 1'b0,  8'd72,  9'd267},{  1'b0, 1'b0,  8'd51,  9'd222},{  1'b0, 1'b0,  8'd45,    9'd0},{  1'b0, 1'b0,  8'd31,  9'd321},{  1'b0, 1'b0,  8'd25,   9'd18},{  1'b0, 1'b0,  8'd15,    9'd0},{  1'b0, 1'b0,  8'd14,   9'd66},{  1'b0, 1'b0,  8'd11,  9'd264},{  1'b0, 1'b0,  8'd10,  9'd332},{  1'b0, 1'b0,   8'd5,  9'd114},{  1'b0, 1'b0,   8'd5,  9'd219},{  1'b0, 1'b1,   8'd0,  9'd213},
{  1'b0, 1'b0, 8'd166,    9'd0},{  1'b0, 1'b0, 8'd165,    9'd0},{  1'b0, 1'b0, 8'd138,  9'd216},{  1'b0, 1'b0, 8'd136,    9'd0},{  1'b0, 1'b0, 8'd129,  9'd211},{  1'b0, 1'b0, 8'd114,   9'd21},{  1'b0, 1'b0, 8'd108,   9'd50},{  1'b0, 1'b0, 8'd106,    9'd0},{  1'b0, 1'b0,  8'd82,  9'd307},{  1'b0, 1'b0,  8'd76,    9'd0},{  1'b0, 1'b0,  8'd61,  9'd112},{  1'b0, 1'b0,  8'd46,    9'd0},{  1'b0, 1'b0,  8'd43,   9'd30},{  1'b0, 1'b0,  8'd36,  9'd348},{  1'b0, 1'b0,  8'd29,  9'd107},{  1'b0, 1'b0,  8'd16,    9'd0},{  1'b0, 1'b0,  8'd14,  9'd181},{  1'b0, 1'b0,   8'd8,  9'd216},{  1'b0, 1'b0,   8'd5,   9'd62},{  1'b0, 1'b0,   8'd2,  9'd290},{  1'b0, 1'b0,   8'd1,   9'd59},{  1'b0, 1'b1,   8'd0,  9'd138},
{  1'b0, 1'b0, 8'd167,    9'd0},{  1'b0, 1'b0, 8'd166,    9'd0},{  1'b0, 1'b0, 8'd149,  9'd267},{  1'b0, 1'b0, 8'd139,  9'd293},{  1'b0, 1'b0, 8'd137,    9'd0},{  1'b0, 1'b0, 8'd107,    9'd0},{  1'b0, 1'b0,  8'd99,  9'd248},{  1'b0, 1'b0,  8'd95,   9'd20},{  1'b0, 1'b0,  8'd77,    9'd0},{  1'b0, 1'b0,  8'd74,  9'd235},{  1'b0, 1'b0,  8'd69,  9'd183},{  1'b0, 1'b0,  8'd47,    9'd0},{  1'b0, 1'b0,  8'd40,  9'd169},{  1'b0, 1'b0,  8'd38,  9'd334},{  1'b0, 1'b0,  8'd26,  9'd127},{  1'b0, 1'b0,  8'd17,    9'd0},{  1'b0, 1'b0,   8'd9,  9'd168},{  1'b0, 1'b0,   8'd6,  9'd130},{  1'b0, 1'b0,   8'd4,   9'd77},{  1'b0, 1'b0,   8'd2,   9'd92},{  1'b0, 1'b0,   8'd1,   9'd98},{  1'b0, 1'b1,   8'd1,  9'd340},
{  1'b0, 1'b0, 8'd168,    9'd0},{  1'b0, 1'b0, 8'd167,    9'd0},{  1'b0, 1'b0, 8'd138,    9'd0},{  1'b0, 1'b0, 8'd134,  9'd305},{  1'b0, 1'b0, 8'd123,  9'd330},{  1'b0, 1'b0, 8'd119,  9'd234},{  1'b0, 1'b0, 8'd108,    9'd0},{  1'b0, 1'b0, 8'd105,   9'd75},{  1'b0, 1'b0,  8'd80,  9'd233},{  1'b0, 1'b0,  8'd78,    9'd0},{  1'b0, 1'b0,  8'd67,  9'd262},{  1'b0, 1'b0,  8'd48,    9'd0},{  1'b0, 1'b0,  8'd41,   9'd28},{  1'b0, 1'b0,  8'd38,  9'd134},{  1'b0, 1'b0,  8'd18,    9'd0},{  1'b0, 1'b0,  8'd16,  9'd216},{  1'b0, 1'b0,  8'd14,   9'd25},{  1'b0, 1'b0,  8'd11,  9'd332},{  1'b0, 1'b0,  8'd10,   9'd61},{  1'b0, 1'b0,   8'd7,  9'd129},{  1'b0, 1'b0,   8'd5,   9'd11},{  1'b0, 1'b1,   8'd3,   9'd37},
{  1'b0, 1'b0, 8'd169,    9'd0},{  1'b0, 1'b0, 8'd168,    9'd0},{  1'b0, 1'b0, 8'd140,   9'd66},{  1'b0, 1'b0, 8'd139,    9'd0},{  1'b0, 1'b0, 8'd122,   9'd78},{  1'b0, 1'b0, 8'd109,    9'd0},{  1'b0, 1'b0, 8'd106,   9'd80},{  1'b0, 1'b0,  8'd94,   9'd64},{  1'b0, 1'b0,  8'd79,    9'd0},{  1'b0, 1'b0,  8'd66,   9'd47},{  1'b0, 1'b0,  8'd60,  9'd118},{  1'b0, 1'b0,  8'd57,  9'd170},{  1'b0, 1'b0,  8'd51,  9'd135},{  1'b0, 1'b0,  8'd49,    9'd0},{  1'b0, 1'b0,  8'd23,  9'd311},{  1'b0, 1'b0,  8'd19,    9'd0},{  1'b0, 1'b0,  8'd10,  9'd212},{  1'b0, 1'b0,   8'd7,  9'd333},{  1'b0, 1'b0,   8'd2,  9'd329},{  1'b0, 1'b0,   8'd1,   9'd82},{  1'b0, 1'b0,   8'd1,  9'd144},{  1'b0, 1'b1,   8'd0,  9'd165},
{  1'b0, 1'b0, 8'd170,    9'd0},{  1'b0, 1'b0, 8'd169,    9'd0},{  1'b0, 1'b0, 8'd140,    9'd0},{  1'b0, 1'b0, 8'd124,  9'd230},{  1'b0, 1'b0, 8'd122,  9'd335},{  1'b0, 1'b0, 8'd110,    9'd0},{  1'b0, 1'b0, 8'd104,  9'd309},{  1'b0, 1'b0,  8'd99,  9'd105},{  1'b0, 1'b0,  8'd80,    9'd0},{  1'b0, 1'b0,  8'd73,  9'd187},{  1'b0, 1'b0,  8'd65,  9'd176},{  1'b0, 1'b0,  8'd50,    9'd0},{  1'b0, 1'b0,  8'd35,   9'd61},{  1'b0, 1'b0,  8'd30,   9'd80},{  1'b0, 1'b0,  8'd26,  9'd286},{  1'b0, 1'b0,  8'd21,   9'd39},{  1'b0, 1'b0,  8'd20,    9'd0},{  1'b0, 1'b0,  8'd14,    9'd6},{  1'b0, 1'b0,   8'd8,  9'd180},{  1'b0, 1'b0,   8'd5,  9'd344},{  1'b0, 1'b0,   8'd5,  9'd195},{  1'b0, 1'b1,   8'd5,   9'd92},
{  1'b0, 1'b0, 8'd171,    9'd0},{  1'b0, 1'b0, 8'd170,    9'd0},{  1'b0, 1'b0, 8'd141,    9'd0},{  1'b0, 1'b0, 8'd126,  9'd260},{  1'b0, 1'b0, 8'd121,  9'd126},{  1'b0, 1'b0, 8'd112,  9'd209},{  1'b0, 1'b0, 8'd111,    9'd0},{  1'b0, 1'b0, 8'd103,  9'd319},{  1'b0, 1'b0,  8'd81,    9'd0},{  1'b0, 1'b0,  8'd70,  9'd164},{  1'b0, 1'b0,  8'd64,   9'd40},{  1'b0, 1'b0,  8'd51,    9'd0},{  1'b0, 1'b0,  8'd33,  9'd177},{  1'b0, 1'b0,  8'd33,   9'd67},{  1'b0, 1'b0,  8'd23,   9'd72},{  1'b0, 1'b0,  8'd21,    9'd0},{  1'b0, 1'b0,  8'd14,  9'd225},{  1'b0, 1'b0,   8'd9,  9'd110},{  1'b0, 1'b0,   8'd8,    9'd3},{  1'b0, 1'b0,   8'd6,  9'd103},{  1'b0, 1'b0,   8'd6,   9'd53},{  1'b0, 1'b1,   8'd4,  9'd243},
{  1'b0, 1'b0, 8'd172,    9'd0},{  1'b0, 1'b0, 8'd171,    9'd0},{  1'b0, 1'b0, 8'd142,    9'd0},{  1'b0, 1'b0, 8'd141,  9'd306},{  1'b0, 1'b0, 8'd134,  9'd303},{  1'b0, 1'b0, 8'd112,    9'd0},{  1'b0, 1'b0, 8'd109,  9'd268},{  1'b0, 1'b0, 8'd101,  9'd357},{  1'b0, 1'b0,  8'd85,  9'd185},{  1'b0, 1'b0,  8'd82,    9'd0},{  1'b0, 1'b0,  8'd81,   9'd53},{  1'b0, 1'b0,  8'd52,    9'd0},{  1'b0, 1'b0,  8'd47,  9'd339},{  1'b0, 1'b0,  8'd32,   9'd81},{  1'b0, 1'b0,  8'd22,    9'd0},{  1'b0, 1'b0,  8'd14,  9'd296},{  1'b0, 1'b0,  8'd13,   9'd82},{  1'b0, 1'b0,  8'd13,   9'd69},{  1'b0, 1'b0,  8'd10,  9'd345},{  1'b0, 1'b0,   8'd9,  9'd329},{  1'b0, 1'b0,   8'd3,  9'd301},{  1'b0, 1'b1,   8'd0,  9'd103},
{  1'b0, 1'b0, 8'd173,    9'd0},{  1'b0, 1'b0, 8'd172,    9'd0},{  1'b0, 1'b0, 8'd143,    9'd0},{  1'b0, 1'b0, 8'd143,  9'd300},{  1'b0, 1'b0, 8'd135,  9'd206},{  1'b0, 1'b0, 8'd114,   9'd76},{  1'b0, 1'b0, 8'd113,    9'd0},{  1'b0, 1'b0, 8'd112,  9'd127},{  1'b0, 1'b0,  8'd84,  9'd124},{  1'b0, 1'b0,  8'd83,    9'd0},{  1'b0, 1'b0,  8'd79,  9'd181},{  1'b0, 1'b0,  8'd54,  9'd282},{  1'b0, 1'b0,  8'd53,    9'd0},{  1'b0, 1'b0,  8'd41,  9'd115},{  1'b0, 1'b0,  8'd23,    9'd0},{  1'b0, 1'b0,  8'd21,  9'd325},{  1'b0, 1'b0,  8'd19,   9'd59},{  1'b0, 1'b0,  8'd14,   9'd36},{  1'b0, 1'b0,  8'd13,  9'd166},{  1'b0, 1'b0,  8'd13,  9'd306},{  1'b0, 1'b0,  8'd10,  9'd243},{  1'b0, 1'b1,   8'd8,  9'd200},
{  1'b0, 1'b0, 8'd174,    9'd0},{  1'b0, 1'b0, 8'd173,    9'd0},{  1'b0, 1'b0, 8'd144,    9'd0},{  1'b0, 1'b0, 8'd142,   9'd57},{  1'b0, 1'b0, 8'd124,   9'd63},{  1'b0, 1'b0, 8'd114,    9'd0},{  1'b0, 1'b0,  8'd96,  9'd284},{  1'b0, 1'b0,  8'd96,   9'd45},{  1'b0, 1'b0,  8'd84,    9'd0},{  1'b0, 1'b0,  8'd68,  9'd342},{  1'b0, 1'b0,  8'd60,   9'd48},{  1'b0, 1'b0,  8'd57,  9'd205},{  1'b0, 1'b0,  8'd54,    9'd0},{  1'b0, 1'b0,  8'd36,  9'd325},{  1'b0, 1'b0,  8'd24,    9'd0},{  1'b0, 1'b0,  8'd20,  9'd205},{  1'b0, 1'b0,  8'd20,  9'd261},{  1'b0, 1'b0,   8'd7,  9'd153},{  1'b0, 1'b0,   8'd4,   9'd26},{  1'b0, 1'b0,   8'd3,  9'd130},{  1'b0, 1'b0,   8'd2,  9'd295},{  1'b0, 1'b1,   8'd1,  9'd182},
{  1'b0, 1'b0, 8'd175,    9'd0},{  1'b0, 1'b0, 8'd174,    9'd0},{  1'b0, 1'b0, 8'd145,    9'd0},{  1'b0, 1'b0, 8'd145,  9'd129},{  1'b0, 1'b0, 8'd139,  9'd254},{  1'b0, 1'b0, 8'd118,   9'd68},{  1'b0, 1'b0, 8'd115,    9'd0},{  1'b0, 1'b0, 8'd110,   9'd69},{  1'b0, 1'b0,  8'd85,    9'd0},{  1'b0, 1'b0,  8'd75,  9'd113},{  1'b0, 1'b0,  8'd68,  9'd147},{  1'b0, 1'b0,  8'd55,    9'd0},{  1'b0, 1'b0,  8'd53,  9'd102},{  1'b0, 1'b0,  8'd30,  9'd234},{  1'b0, 1'b0,  8'd25,    9'd0},{  1'b0, 1'b0,  8'd13,  9'd336},{  1'b0, 1'b0,  8'd12,  9'd259},{  1'b0, 1'b0,  8'd12,  9'd303},{  1'b0, 1'b0,  8'd11,   9'd79},{  1'b0, 1'b0,  8'd10,  9'd152},{  1'b0, 1'b0,   8'd3,  9'd159},{  1'b0, 1'b1,   8'd3,  9'd338},
{  1'b0, 1'b0, 8'd176,    9'd0},{  1'b0, 1'b0, 8'd175,    9'd0},{  1'b0, 1'b0, 8'd147,  9'd317},{  1'b0, 1'b0, 8'd146,    9'd0},{  1'b0, 1'b0, 8'd138,  9'd351},{  1'b0, 1'b0, 8'd116,    9'd0},{  1'b0, 1'b0,  8'd97,  9'd355},{  1'b0, 1'b0,  8'd95,    9'd6},{  1'b0, 1'b0,  8'd86,    9'd0},{  1'b0, 1'b0,  8'd78,  9'd206},{  1'b0, 1'b0,  8'd76,  9'd128},{  1'b0, 1'b0,  8'd56,    9'd0},{  1'b0, 1'b0,  8'd52,   9'd33},{  1'b0, 1'b0,  8'd50,  9'd158},{  1'b0, 1'b0,  8'd26,    9'd0},{  1'b0, 1'b0,  8'd25,   9'd51},{  1'b0, 1'b0,  8'd10,  9'd217},{  1'b0, 1'b0,  8'd10,   9'd58},{  1'b0, 1'b0,  8'd10,   9'd81},{  1'b0, 1'b0,  8'd10,  9'd186},{  1'b0, 1'b0,   8'd6,  9'd115},{  1'b0, 1'b1,   8'd0,   9'd13},
{  1'b0, 1'b0, 8'd177,    9'd0},{  1'b0, 1'b0, 8'd176,    9'd0},{  1'b0, 1'b0, 8'd149,  9'd244},{  1'b0, 1'b0, 8'd147,    9'd0},{  1'b0, 1'b0, 8'd131,  9'd260},{  1'b0, 1'b0, 8'd117,    9'd0},{  1'b0, 1'b0, 8'd107,   9'd51},{  1'b0, 1'b0, 8'd104,  9'd208},{  1'b0, 1'b0,  8'd87,    9'd0},{  1'b0, 1'b0,  8'd84,  9'd307},{  1'b0, 1'b0,  8'd75,  9'd300},{  1'b0, 1'b0,  8'd57,    9'd0},{  1'b0, 1'b0,  8'd50,   9'd89},{  1'b0, 1'b0,  8'd44,  9'd136},{  1'b0, 1'b0,  8'd27,    9'd0},{  1'b0, 1'b0,  8'd14,  9'd150},{  1'b0, 1'b0,  8'd12,  9'd228},{  1'b0, 1'b0,  8'd12,  9'd213},{  1'b0, 1'b0,  8'd11,  9'd308},{  1'b0, 1'b0,   8'd8,  9'd352},{  1'b0, 1'b0,   8'd7,  9'd107},{  1'b0, 1'b1,   8'd4,  9'd238},
{  1'b0, 1'b0, 8'd178,    9'd0},{  1'b0, 1'b0, 8'd177,    9'd0},{  1'b0, 1'b0, 8'd148,    9'd0},{  1'b0, 1'b0, 8'd128,  9'd182},{  1'b0, 1'b0, 8'd127,  9'd254},{  1'b0, 1'b0, 8'd118,    9'd0},{  1'b0, 1'b0, 8'd110,  9'd298},{  1'b0, 1'b0,  8'd92,   9'd10},{  1'b0, 1'b0,  8'd88,    9'd0},{  1'b0, 1'b0,  8'd85,  9'd233},{  1'b0, 1'b0,  8'd74,  9'd295},{  1'b0, 1'b0,  8'd58,    9'd0},{  1'b0, 1'b0,  8'd48,  9'd188},{  1'b0, 1'b0,  8'd35,   9'd77},{  1'b0, 1'b0,  8'd28,    9'd0},{  1'b0, 1'b0,  8'd18,   9'd56},{  1'b0, 1'b0,  8'd14,  9'd323},{  1'b0, 1'b0,  8'd11,  9'd198},{  1'b0, 1'b0,  8'd10,  9'd284},{  1'b0, 1'b0,   8'd8,   9'd98},{  1'b0, 1'b0,   8'd4,   9'd50},{  1'b0, 1'b1,   8'd1,  9'd242},
{  1'b0, 1'b0, 8'd179,    9'd0},{  1'b0, 1'b0, 8'd178,    9'd0},{  1'b0, 1'b0, 8'd149,    9'd0},{  1'b0, 1'b0, 8'd125,  9'd188},{  1'b0, 1'b0, 8'd120,   9'd58},{  1'b0, 1'b0, 8'd119,    9'd0},{  1'b0, 1'b0,  8'd93,   9'd73},{  1'b0, 1'b0,  8'd93,  9'd309},{  1'b0, 1'b0,  8'd89,    9'd0},{  1'b0, 1'b0,  8'd88,  9'd268},{  1'b0, 1'b0,  8'd66,  9'd324},{  1'b0, 1'b0,  8'd59,    9'd0},{  1'b0, 1'b0,  8'd49,  9'd114},{  1'b0, 1'b0,  8'd44,   9'd51},{  1'b0, 1'b0,  8'd29,    9'd0},{  1'b0, 1'b0,  8'd24,   9'd64},{  1'b0, 1'b0,  8'd16,  9'd306},{  1'b0, 1'b0,  8'd11,  9'd242},{  1'b0, 1'b0,   8'd6,  9'd197},{  1'b0, 1'b0,   8'd4,   9'd10},{  1'b0, 1'b0,   8'd2,   9'd72},{  1'b0, 1'b1,   8'd0,  9'd296}
};
localparam bit [18 : 0] cLARGE_HS_V_TAB_5BY6_PACKED[cLARGE_HS_TAB_5BY6_PACKED_SIZE] = '{
{8'd179, 1'b0,   10'd0},{8'd179, 1'b1, 10'd638},
{8'd178, 1'b0, 10'd616},{8'd178, 1'b1, 10'd639},
{8'd177, 1'b0, 10'd594},{8'd177, 1'b1, 10'd617},
{8'd176, 1'b0, 10'd572},{8'd176, 1'b1, 10'd595},
{8'd175, 1'b0, 10'd550},{8'd175, 1'b1, 10'd573},
{8'd174, 1'b0, 10'd528},{8'd174, 1'b1, 10'd551},
{8'd173, 1'b0, 10'd506},{8'd173, 1'b1, 10'd529},
{8'd172, 1'b0, 10'd484},{8'd172, 1'b1, 10'd507},
{8'd171, 1'b0, 10'd462},{8'd171, 1'b1, 10'd485},
{8'd170, 1'b0, 10'd440},{8'd170, 1'b1, 10'd463},
{8'd169, 1'b0, 10'd418},{8'd169, 1'b1, 10'd441},
{8'd168, 1'b0, 10'd396},{8'd168, 1'b1, 10'd419},
{8'd167, 1'b0, 10'd374},{8'd167, 1'b1, 10'd397},
{8'd166, 1'b0, 10'd352},{8'd166, 1'b1, 10'd375},
{8'd165, 1'b0, 10'd330},{8'd165, 1'b1, 10'd353},
{8'd164, 1'b0, 10'd308},{8'd164, 1'b1, 10'd331},
{8'd163, 1'b0, 10'd286},{8'd163, 1'b1, 10'd309},
{8'd162, 1'b0, 10'd264},{8'd162, 1'b1, 10'd287},
{8'd161, 1'b0, 10'd242},{8'd161, 1'b1, 10'd265},
{8'd160, 1'b0, 10'd220},{8'd160, 1'b1, 10'd243},
{8'd159, 1'b0, 10'd198},{8'd159, 1'b1, 10'd221},
{8'd158, 1'b0, 10'd176},{8'd158, 1'b1, 10'd199},
{8'd157, 1'b0, 10'd154},{8'd157, 1'b1, 10'd177},
{8'd156, 1'b0, 10'd132},{8'd156, 1'b1, 10'd155},
{8'd155, 1'b0, 10'd110},{8'd155, 1'b1, 10'd133},
{8'd154, 1'b0,  10'd88},{8'd154, 1'b1, 10'd111},
{8'd153, 1'b0,  10'd66},{8'd153, 1'b1,  10'd89},
{8'd152, 1'b0,  10'd44},{8'd152, 1'b1,  10'd67},
{8'd151, 1'b0,  10'd22},{8'd151, 1'b1,  10'd45},
{8'd150, 1'b0,   10'd1},{8'd150, 1'b1,  10'd23},
{8'd149, 1'b0, 10'd376},{8'd149, 1'b0, 10'd596},{8'd149, 1'b1, 10'd640},
{8'd148, 1'b0,  10'd24},{8'd148, 1'b0,  10'd68},{8'd148, 1'b1, 10'd618},
{8'd147, 1'b0, 10'd112},{8'd147, 1'b0, 10'd574},{8'd147, 1'b1, 10'd597},
{8'd146, 1'b0,  10'd90},{8'd146, 1'b0, 10'd266},{8'd146, 1'b1, 10'd575},
{8'd145, 1'b0, 10'd244},{8'd145, 1'b0, 10'd552},{8'd145, 1'b1, 10'd553},
{8'd144, 1'b0, 10'd245},{8'd144, 1'b0, 10'd288},{8'd144, 1'b1, 10'd530},
{8'd143, 1'b0, 10'd134},{8'd143, 1'b0, 10'd508},{8'd143, 1'b1, 10'd509},
{8'd142, 1'b0, 10'd289},{8'd142, 1'b0, 10'd486},{8'd142, 1'b1, 10'd531},
{8'd141, 1'b0, 10'd178},{8'd141, 1'b0, 10'd464},{8'd141, 1'b1, 10'd487},
{8'd140, 1'b0,   10'd2},{8'd140, 1'b0, 10'd420},{8'd140, 1'b1, 10'd442},
{8'd139, 1'b0, 10'd377},{8'd139, 1'b0, 10'd421},{8'd139, 1'b1, 10'd554},
{8'd138, 1'b0, 10'd354},{8'd138, 1'b0, 10'd398},{8'd138, 1'b1, 10'd576},
{8'd137, 1'b0,  10'd69},{8'd137, 1'b0,  10'd91},{8'd137, 1'b1, 10'd378},
{8'd136, 1'b0,   10'd3},{8'd136, 1'b0, 10'd332},{8'd136, 1'b1, 10'd355},
{8'd135, 1'b0, 10'd267},{8'd135, 1'b0, 10'd333},{8'd135, 1'b1, 10'd510},
{8'd134, 1'b0, 10'd310},{8'd134, 1'b0, 10'd399},{8'd134, 1'b1, 10'd488},
{8'd133, 1'b0, 10'd200},{8'd133, 1'b0, 10'd222},{8'd133, 1'b1, 10'd290},
{8'd132, 1'b0,  10'd46},{8'd132, 1'b0, 10'd113},{8'd132, 1'b1, 10'd268},
{8'd131, 1'b0,  10'd25},{8'd131, 1'b0, 10'd246},{8'd131, 1'b1, 10'd598},
{8'd130, 1'b0,  10'd47},{8'd130, 1'b0, 10'd179},{8'd130, 1'b1, 10'd223},
{8'd129, 1'b0, 10'd135},{8'd129, 1'b0, 10'd201},{8'd129, 1'b1, 10'd356},
{8'd128, 1'b0, 10'd180},{8'd128, 1'b0, 10'd224},{8'd128, 1'b1, 10'd619},
{8'd127, 1'b0, 10'd156},{8'd127, 1'b0, 10'd311},{8'd127, 1'b1, 10'd620},
{8'd126, 1'b0, 10'd136},{8'd126, 1'b0, 10'd334},{8'd126, 1'b1, 10'd465},
{8'd125, 1'b0, 10'd114},{8'd125, 1'b0, 10'd312},{8'd125, 1'b1, 10'd641},
{8'd124, 1'b0,  10'd92},{8'd124, 1'b0, 10'd443},{8'd124, 1'b1, 10'd532},
{8'd123, 1'b0,  10'd70},{8'd123, 1'b0, 10'd157},{8'd123, 1'b1, 10'd400},
{8'd122, 1'b0,  10'd48},{8'd122, 1'b0, 10'd422},{8'd122, 1'b1, 10'd444},
{8'd121, 1'b0,  10'd26},{8'd121, 1'b0, 10'd202},{8'd121, 1'b1, 10'd466},
{8'd120, 1'b0,   10'd4},{8'd120, 1'b0, 10'd158},{8'd120, 1'b1, 10'd642},
{8'd119, 1'b0, 10'd291},{8'd119, 1'b0, 10'd401},{8'd119, 1'b1, 10'd643},
{8'd118, 1'b0,   10'd5},{8'd118, 1'b0, 10'd555},{8'd118, 1'b1, 10'd621},
{8'd117, 1'b0, 10'd225},{8'd117, 1'b0, 10'd313},{8'd117, 1'b1, 10'd599},
{8'd116, 1'b0,  10'd49},{8'd116, 1'b0, 10'd159},{8'd116, 1'b1, 10'd577},
{8'd115, 1'b0, 10'd115},{8'd115, 1'b0, 10'd247},{8'd115, 1'b1, 10'd556},
{8'd114, 1'b0, 10'd357},{8'd114, 1'b0, 10'd511},{8'd114, 1'b1, 10'd533},
{8'd113, 1'b0,  10'd93},{8'd113, 1'b0, 10'd314},{8'd113, 1'b1, 10'd512},
{8'd112, 1'b0, 10'd467},{8'd112, 1'b0, 10'd489},{8'd112, 1'b1, 10'd513},
{8'd111, 1'b0,  10'd71},{8'd111, 1'b0, 10'd137},{8'd111, 1'b1, 10'd468},
{8'd110, 1'b0, 10'd445},{8'd110, 1'b0, 10'd557},{8'd110, 1'b1, 10'd622},
{8'd109, 1'b0,  10'd94},{8'd109, 1'b0, 10'd423},{8'd109, 1'b1, 10'd490},
{8'd108, 1'b0, 10'd335},{8'd108, 1'b0, 10'd358},{8'd108, 1'b1, 10'd402},
{8'd107, 1'b0, 10'd138},{8'd107, 1'b0, 10'd379},{8'd107, 1'b1, 10'd600},
{8'd106, 1'b0, 10'd336},{8'd106, 1'b0, 10'd359},{8'd106, 1'b1, 10'd424},
{8'd105, 1'b0, 10'd203},{8'd105, 1'b0, 10'd337},{8'd105, 1'b1, 10'd403},
{8'd104, 1'b0, 10'd315},{8'd104, 1'b0, 10'd446},{8'd104, 1'b1, 10'd601},
{8'd103, 1'b0, 10'd226},{8'd103, 1'b0, 10'd292},{8'd103, 1'b1, 10'd469},
{8'd102, 1'b0, 10'd269},{8'd102, 1'b0, 10'd270},{8'd102, 1'b1, 10'd293},
{8'd101, 1'b0,  10'd27},{8'd101, 1'b0, 10'd248},{8'd101, 1'b1, 10'd491},
{8'd100, 1'b0,  10'd28},{8'd100, 1'b0, 10'd181},{8'd100, 1'b1, 10'd227},
{ 8'd99, 1'b0, 10'd204},{ 8'd99, 1'b0, 10'd380},{ 8'd99, 1'b1, 10'd447},
{ 8'd98, 1'b0, 10'd182},{ 8'd98, 1'b0, 10'd205},{ 8'd98, 1'b1, 10'd271},
{ 8'd97, 1'b0,   10'd6},{ 8'd97, 1'b0, 10'd160},{ 8'd97, 1'b1, 10'd578},
{ 8'd96, 1'b0, 10'd139},{ 8'd96, 1'b0, 10'd534},{ 8'd96, 1'b1, 10'd535},
{ 8'd95, 1'b0, 10'd116},{ 8'd95, 1'b0, 10'd381},{ 8'd95, 1'b1, 10'd579},
{ 8'd94, 1'b0,  10'd95},{ 8'd94, 1'b0, 10'd183},{ 8'd94, 1'b1, 10'd425},
{ 8'd93, 1'b0,  10'd72},{ 8'd93, 1'b0, 10'd644},{ 8'd93, 1'b1, 10'd645},
{ 8'd92, 1'b0,  10'd50},{ 8'd92, 1'b0, 10'd161},{ 8'd92, 1'b1, 10'd623},
{ 8'd91, 1'b0,  10'd29},{ 8'd91, 1'b0,  10'd51},{ 8'd91, 1'b1, 10'd117},
{ 8'd90, 1'b0,   10'd7},{ 8'd90, 1'b0,  10'd73},{ 8'd90, 1'b1, 10'd249},
{ 8'd89, 1'b0, 10'd118},{ 8'd89, 1'b0, 10'd250},{ 8'd89, 1'b1, 10'd646},
{ 8'd88, 1'b0, 10'd294},{ 8'd88, 1'b0, 10'd624},{ 8'd88, 1'b1, 10'd647},
{ 8'd87, 1'b0,  10'd96},{ 8'd87, 1'b0, 10'd295},{ 8'd87, 1'b1, 10'd602},
{ 8'd86, 1'b0, 10'd140},{ 8'd86, 1'b0, 10'd272},{ 8'd86, 1'b1, 10'd580},
{ 8'd85, 1'b0, 10'd492},{ 8'd85, 1'b0, 10'd558},{ 8'd85, 1'b1, 10'd625},
{ 8'd84, 1'b0, 10'd514},{ 8'd84, 1'b0, 10'd536},{ 8'd84, 1'b1, 10'd603},
{ 8'd83, 1'b0, 10'd162},{ 8'd83, 1'b0, 10'd228},{ 8'd83, 1'b1, 10'd515},
{ 8'd82, 1'b0, 10'd206},{ 8'd82, 1'b0, 10'd360},{ 8'd82, 1'b1, 10'd493},
{ 8'd81, 1'b0, 10'd273},{ 8'd81, 1'b0, 10'd470},{ 8'd81, 1'b1, 10'd494},
{ 8'd80, 1'b0, 10'd338},{ 8'd80, 1'b0, 10'd404},{ 8'd80, 1'b1, 10'd448},
{ 8'd79, 1'b0,  10'd74},{ 8'd79, 1'b0, 10'd426},{ 8'd79, 1'b1, 10'd516},
{ 8'd78, 1'b0,   10'd8},{ 8'd78, 1'b0, 10'd405},{ 8'd78, 1'b1, 10'd581},
{ 8'd77, 1'b0,  10'd97},{ 8'd77, 1'b0, 10'd207},{ 8'd77, 1'b1, 10'd382},
{ 8'd76, 1'b0, 10'd229},{ 8'd76, 1'b0, 10'd361},{ 8'd76, 1'b1, 10'd582},
{ 8'd75, 1'b0, 10'd339},{ 8'd75, 1'b0, 10'd559},{ 8'd75, 1'b1, 10'd604},
{ 8'd74, 1'b0, 10'd316},{ 8'd74, 1'b0, 10'd383},{ 8'd74, 1'b1, 10'd626},
{ 8'd73, 1'b0, 10'd141},{ 8'd73, 1'b0, 10'd296},{ 8'd73, 1'b1, 10'd449},
{ 8'd72, 1'b0,   10'd9},{ 8'd72, 1'b0, 10'd274},{ 8'd72, 1'b1, 10'd340},
{ 8'd71, 1'b0, 10'd184},{ 8'd71, 1'b0, 10'd251},{ 8'd71, 1'b1, 10'd317},
{ 8'd70, 1'b0,  10'd52},{ 8'd70, 1'b0, 10'd230},{ 8'd70, 1'b1, 10'd471},
{ 8'd69, 1'b0,  10'd30},{ 8'd69, 1'b0, 10'd208},{ 8'd69, 1'b1, 10'd384},
{ 8'd68, 1'b0, 10'd185},{ 8'd68, 1'b0, 10'd537},{ 8'd68, 1'b1, 10'd560},
{ 8'd67, 1'b0,  10'd31},{ 8'd67, 1'b0, 10'd163},{ 8'd67, 1'b1, 10'd406},
{ 8'd66, 1'b0, 10'd142},{ 8'd66, 1'b0, 10'd427},{ 8'd66, 1'b1, 10'd648},
{ 8'd65, 1'b0,  10'd53},{ 8'd65, 1'b0, 10'd119},{ 8'd65, 1'b1, 10'd450},
{ 8'd64, 1'b0,  10'd75},{ 8'd64, 1'b0,  10'd98},{ 8'd64, 1'b1, 10'd472},
{ 8'd63, 1'b0,  10'd76},{ 8'd63, 1'b0, 10'd120},{ 8'd63, 1'b1, 10'd252},
{ 8'd62, 1'b0,  10'd54},{ 8'd62, 1'b0, 10'd164},{ 8'd62, 1'b1, 10'd186},
{ 8'd61, 1'b0,  10'd32},{ 8'd61, 1'b0, 10'd318},{ 8'd61, 1'b1, 10'd362},
{ 8'd60, 1'b0,  10'd10},{ 8'd60, 1'b0, 10'd428},{ 8'd60, 1'b1, 10'd538},
{ 8'd59, 1'b0, 10'd253},{ 8'd59, 1'b0, 10'd319},{ 8'd59, 1'b1, 10'd649},
{ 8'd58, 1'b0,  10'd77},{ 8'd58, 1'b0, 10'd209},{ 8'd58, 1'b1, 10'd627},
{ 8'd57, 1'b0, 10'd429},{ 8'd57, 1'b0, 10'd539},{ 8'd57, 1'b1, 10'd605},
{ 8'd56, 1'b0,  10'd55},{ 8'd56, 1'b0, 10'd187},{ 8'd56, 1'b1, 10'd583},
{ 8'd55, 1'b0,  10'd99},{ 8'd55, 1'b0, 10'd121},{ 8'd55, 1'b1, 10'd561},
{ 8'd54, 1'b0,  10'd11},{ 8'd54, 1'b0, 10'd517},{ 8'd54, 1'b1, 10'd540},
{ 8'd53, 1'b0, 10'd210},{ 8'd53, 1'b0, 10'd518},{ 8'd53, 1'b1, 10'd562},
{ 8'd52, 1'b0, 10'd165},{ 8'd52, 1'b0, 10'd495},{ 8'd52, 1'b1, 10'd584},
{ 8'd51, 1'b0, 10'd341},{ 8'd51, 1'b0, 10'd430},{ 8'd51, 1'b1, 10'd473},
{ 8'd50, 1'b0, 10'd451},{ 8'd50, 1'b0, 10'd585},{ 8'd50, 1'b1, 10'd606},
{ 8'd49, 1'b0, 10'd231},{ 8'd49, 1'b0, 10'd431},{ 8'd49, 1'b1, 10'd650},
{ 8'd48, 1'b0, 10'd122},{ 8'd48, 1'b0, 10'd407},{ 8'd48, 1'b1, 10'd628},
{ 8'd47, 1'b0, 10'd166},{ 8'd47, 1'b0, 10'd385},{ 8'd47, 1'b1, 10'd496},
{ 8'd46, 1'b0,  10'd33},{ 8'd46, 1'b0, 10'd275},{ 8'd46, 1'b1, 10'd363},
{ 8'd45, 1'b0, 10'd143},{ 8'd45, 1'b0, 10'd254},{ 8'd45, 1'b1, 10'd342},
{ 8'd44, 1'b0, 10'd320},{ 8'd44, 1'b0, 10'd607},{ 8'd44, 1'b1, 10'd651},
{ 8'd43, 1'b0, 10'd297},{ 8'd43, 1'b0, 10'd298},{ 8'd43, 1'b1, 10'd364},
{ 8'd42, 1'b0,  10'd56},{ 8'd42, 1'b0, 10'd276},{ 8'd42, 1'b1, 10'd299},
{ 8'd41, 1'b0, 10'd255},{ 8'd41, 1'b0, 10'd408},{ 8'd41, 1'b1, 10'd519},
{ 8'd40, 1'b0,  10'd12},{ 8'd40, 1'b0, 10'd232},{ 8'd40, 1'b1, 10'd386},
{ 8'd39, 1'b0, 10'd100},{ 8'd39, 1'b0, 10'd188},{ 8'd39, 1'b1, 10'd211},
{ 8'd38, 1'b0, 10'd189},{ 8'd38, 1'b0, 10'd387},{ 8'd38, 1'b1, 10'd409},
{ 8'd37, 1'b0, 10'd144},{ 8'd37, 1'b0, 10'd167},{ 8'd37, 1'b1, 10'd277},
{ 8'd36, 1'b0, 10'd145},{ 8'd36, 1'b0, 10'd365},{ 8'd36, 1'b1, 10'd541},
{ 8'd35, 1'b0, 10'd123},{ 8'd35, 1'b0, 10'd452},{ 8'd35, 1'b1, 10'd629},
{ 8'd34, 1'b0,  10'd78},{ 8'd34, 1'b0, 10'd101},{ 8'd34, 1'b1, 10'd233},
{ 8'd33, 1'b0,  10'd79},{ 8'd33, 1'b0, 10'd474},{ 8'd33, 1'b1, 10'd475},
{ 8'd32, 1'b0,  10'd57},{ 8'd32, 1'b0, 10'd321},{ 8'd32, 1'b1, 10'd497},
{ 8'd31, 1'b0,  10'd34},{ 8'd31, 1'b0,  10'd35},{ 8'd31, 1'b1, 10'd343},
{ 8'd30, 1'b0,  10'd13},{ 8'd30, 1'b0, 10'd453},{ 8'd30, 1'b1, 10'd563},
{ 8'd29, 1'b0, 10'd278},{ 8'd29, 1'b0, 10'd366},{ 8'd29, 1'b1, 10'd652},
{ 8'd28, 1'b0,  10'd58},{ 8'd28, 1'b0, 10'd190},{ 8'd28, 1'b1, 10'd630},
{ 8'd27, 1'b0,  10'd59},{ 8'd27, 1'b0, 10'd168},{ 8'd27, 1'b1, 10'd608},
{ 8'd26, 1'b0, 10'd388},{ 8'd26, 1'b0, 10'd454},{ 8'd26, 1'b1, 10'd586},
{ 8'd25, 1'b0, 10'd344},{ 8'd25, 1'b0, 10'd564},{ 8'd25, 1'b1, 10'd587},
{ 8'd24, 1'b0, 10'd234},{ 8'd24, 1'b0, 10'd542},{ 8'd24, 1'b1, 10'd653},
{ 8'd23, 1'b0, 10'd432},{ 8'd23, 1'b0, 10'd476},{ 8'd23, 1'b1, 10'd520},
{ 8'd22, 1'b0, 10'd169},{ 8'd22, 1'b0, 10'd191},{ 8'd22, 1'b1, 10'd498},
{ 8'd21, 1'b0, 10'd455},{ 8'd21, 1'b0, 10'd477},{ 8'd21, 1'b1, 10'd521},
{ 8'd20, 1'b0, 10'd456},{ 8'd20, 1'b0, 10'd543},{ 8'd20, 1'b1, 10'd544},
{ 8'd19, 1'b0,  10'd36},{ 8'd19, 1'b0, 10'd433},{ 8'd19, 1'b1, 10'd522},
{ 8'd18, 1'b0, 10'd235},{ 8'd18, 1'b0, 10'd410},{ 8'd18, 1'b1, 10'd631},
{ 8'd17, 1'b0,  10'd80},{ 8'd17, 1'b0, 10'd146},{ 8'd17, 1'b1, 10'd389},
{ 8'd16, 1'b0, 10'd367},{ 8'd16, 1'b0, 10'd411},{ 8'd16, 1'b1, 10'd654},
{ 8'd15, 1'b0,  10'd37},{ 8'd15, 1'b0, 10'd102},{ 8'd15, 1'b1, 10'd345},
{ 8'd14, 1'b0,  10'd14},{ 8'd14, 1'b0,  10'd15},{ 8'd14, 1'b0, 10'd236},{ 8'd14, 1'b0, 10'd322},{ 8'd14, 1'b0, 10'd346},{ 8'd14, 1'b0, 10'd368},{ 8'd14, 1'b0, 10'd412},{ 8'd14, 1'b0, 10'd457},{ 8'd14, 1'b0, 10'd478},{ 8'd14, 1'b0, 10'd499},{ 8'd14, 1'b0, 10'd523},{ 8'd14, 1'b0, 10'd609},{ 8'd14, 1'b1, 10'd632},
{ 8'd13, 1'b0,  10'd16},{ 8'd13, 1'b0,  10'd38},{ 8'd13, 1'b0, 10'd124},{ 8'd13, 1'b0, 10'd192},{ 8'd13, 1'b0, 10'd212},{ 8'd13, 1'b0, 10'd256},{ 8'd13, 1'b0, 10'd300},{ 8'd13, 1'b0, 10'd301},{ 8'd13, 1'b0, 10'd500},{ 8'd13, 1'b0, 10'd501},{ 8'd13, 1'b0, 10'd524},{ 8'd13, 1'b0, 10'd525},{ 8'd13, 1'b1, 10'd565},
{ 8'd12, 1'b0,  10'd60},{ 8'd12, 1'b0,  10'd61},{ 8'd12, 1'b0,  10'd81},{ 8'd12, 1'b0, 10'd125},{ 8'd12, 1'b0, 10'd193},{ 8'd12, 1'b0, 10'd257},{ 8'd12, 1'b0, 10'd279},{ 8'd12, 1'b0, 10'd302},{ 8'd12, 1'b0, 10'd323},{ 8'd12, 1'b0, 10'd566},{ 8'd12, 1'b0, 10'd567},{ 8'd12, 1'b0, 10'd610},{ 8'd12, 1'b1, 10'd611},
{ 8'd11, 1'b0,  10'd82},{ 8'd11, 1'b0, 10'd103},{ 8'd11, 1'b0, 10'd147},{ 8'd11, 1'b0, 10'd258},{ 8'd11, 1'b0, 10'd259},{ 8'd11, 1'b0, 10'd280},{ 8'd11, 1'b0, 10'd324},{ 8'd11, 1'b0, 10'd347},{ 8'd11, 1'b0, 10'd413},{ 8'd11, 1'b0, 10'd568},{ 8'd11, 1'b0, 10'd612},{ 8'd11, 1'b0, 10'd633},{ 8'd11, 1'b1, 10'd655},
{ 8'd10, 1'b0, 10'd237},{ 8'd10, 1'b0, 10'd281},{ 8'd10, 1'b0, 10'd348},{ 8'd10, 1'b0, 10'd414},{ 8'd10, 1'b0, 10'd434},{ 8'd10, 1'b0, 10'd502},{ 8'd10, 1'b0, 10'd526},{ 8'd10, 1'b0, 10'd569},{ 8'd10, 1'b0, 10'd588},{ 8'd10, 1'b0, 10'd589},{ 8'd10, 1'b0, 10'd590},{ 8'd10, 1'b0, 10'd591},{ 8'd10, 1'b1, 10'd634},
{  8'd9, 1'b0,  10'd17},{  8'd9, 1'b0,  10'd62},{  8'd9, 1'b0, 10'd104},{  8'd9, 1'b0, 10'd105},{  8'd9, 1'b0, 10'd148},{  8'd9, 1'b0, 10'd213},{  8'd9, 1'b0, 10'd238},{  8'd9, 1'b0, 10'd282},{  8'd9, 1'b0, 10'd303},{  8'd9, 1'b0, 10'd325},{  8'd9, 1'b0, 10'd390},{  8'd9, 1'b0, 10'd479},{  8'd9, 1'b1, 10'd503},
{  8'd8, 1'b0,  10'd18},{  8'd8, 1'b0,  10'd83},{  8'd8, 1'b0, 10'd106},{  8'd8, 1'b0, 10'd126},{  8'd8, 1'b0, 10'd194},{  8'd8, 1'b0, 10'd214},{  8'd8, 1'b0, 10'd215},{  8'd8, 1'b0, 10'd369},{  8'd8, 1'b0, 10'd458},{  8'd8, 1'b0, 10'd480},{  8'd8, 1'b0, 10'd527},{  8'd8, 1'b0, 10'd613},{  8'd8, 1'b1, 10'd635},
{  8'd7, 1'b0,  10'd39},{  8'd7, 1'b0, 10'd127},{  8'd7, 1'b0, 10'd149},{  8'd7, 1'b0, 10'd170},{  8'd7, 1'b0, 10'd171},{  8'd7, 1'b0, 10'd172},{  8'd7, 1'b0, 10'd283},{  8'd7, 1'b0, 10'd304},{  8'd7, 1'b0, 10'd326},{  8'd7, 1'b0, 10'd415},{  8'd7, 1'b0, 10'd435},{  8'd7, 1'b0, 10'd545},{  8'd7, 1'b1, 10'd614},
{  8'd6, 1'b0,  10'd19},{  8'd6, 1'b0, 10'd150},{  8'd6, 1'b0, 10'd151},{  8'd6, 1'b0, 10'd216},{  8'd6, 1'b0, 10'd217},{  8'd6, 1'b0, 10'd260},{  8'd6, 1'b0, 10'd261},{  8'd6, 1'b0, 10'd327},{  8'd6, 1'b0, 10'd391},{  8'd6, 1'b0, 10'd481},{  8'd6, 1'b0, 10'd482},{  8'd6, 1'b0, 10'd592},{  8'd6, 1'b1, 10'd656},
{  8'd5, 1'b0,  10'd63},{  8'd5, 1'b0,  10'd84},{  8'd5, 1'b0, 10'd107},{  8'd5, 1'b0, 10'd128},{  8'd5, 1'b0, 10'd262},{  8'd5, 1'b0, 10'd328},{  8'd5, 1'b0, 10'd349},{  8'd5, 1'b0, 10'd350},{  8'd5, 1'b0, 10'd370},{  8'd5, 1'b0, 10'd416},{  8'd5, 1'b0, 10'd459},{  8'd5, 1'b0, 10'd460},{  8'd5, 1'b1, 10'd461},
{  8'd4, 1'b0,  10'd85},{  8'd4, 1'b0, 10'd108},{  8'd4, 1'b0, 10'd109},{  8'd4, 1'b0, 10'd129},{  8'd4, 1'b0, 10'd218},{  8'd4, 1'b0, 10'd239},{  8'd4, 1'b0, 10'd305},{  8'd4, 1'b0, 10'd392},{  8'd4, 1'b0, 10'd483},{  8'd4, 1'b0, 10'd546},{  8'd4, 1'b0, 10'd615},{  8'd4, 1'b0, 10'd636},{  8'd4, 1'b1, 10'd657},
{  8'd3, 1'b0,  10'd20},{  8'd3, 1'b0,  10'd86},{  8'd3, 1'b0, 10'd152},{  8'd3, 1'b0, 10'd173},{  8'd3, 1'b0, 10'd195},{  8'd3, 1'b0, 10'd196},{  8'd3, 1'b0, 10'd240},{  8'd3, 1'b0, 10'd329},{  8'd3, 1'b0, 10'd417},{  8'd3, 1'b0, 10'd504},{  8'd3, 1'b0, 10'd547},{  8'd3, 1'b0, 10'd570},{  8'd3, 1'b1, 10'd571},
{  8'd2, 1'b0,  10'd40},{  8'd2, 1'b0,  10'd41},{  8'd2, 1'b0,  10'd64},{  8'd2, 1'b0, 10'd130},{  8'd2, 1'b0, 10'd131},{  8'd2, 1'b0, 10'd174},{  8'd2, 1'b0, 10'd219},{  8'd2, 1'b0, 10'd284},{  8'd2, 1'b0, 10'd371},{  8'd2, 1'b0, 10'd393},{  8'd2, 1'b0, 10'd436},{  8'd2, 1'b0, 10'd548},{  8'd2, 1'b1, 10'd658},
{  8'd1, 1'b0,  10'd42},{  8'd1, 1'b0,  10'd43},{  8'd1, 1'b0, 10'd175},{  8'd1, 1'b0, 10'd197},{  8'd1, 1'b0, 10'd263},{  8'd1, 1'b0, 10'd306},{  8'd1, 1'b0, 10'd372},{  8'd1, 1'b0, 10'd394},{  8'd1, 1'b0, 10'd395},{  8'd1, 1'b0, 10'd437},{  8'd1, 1'b0, 10'd438},{  8'd1, 1'b0, 10'd549},{  8'd1, 1'b1, 10'd637},
{  8'd0, 1'b0,  10'd21},{  8'd0, 1'b0,  10'd65},{  8'd0, 1'b0,  10'd87},{  8'd0, 1'b0, 10'd153},{  8'd0, 1'b0, 10'd241},{  8'd0, 1'b0, 10'd285},{  8'd0, 1'b0, 10'd307},{  8'd0, 1'b0, 10'd351},{  8'd0, 1'b0, 10'd373},{  8'd0, 1'b0, 10'd439},{  8'd0, 1'b0, 10'd505},{  8'd0, 1'b0, 10'd593},{  8'd0, 1'b1, 10'd659}
};
localparam int          cLARGE_HS_TAB_8BY9_PACKED_SIZE = 540;
localparam bit [18 : 0] cLARGE_HS_TAB_8BY9_PACKED[cLARGE_HS_TAB_8BY9_PACKED_SIZE] = '{
{  1'b1, 1'b0, 8'd179,    9'd1},{  1'b0, 1'b0, 8'd160,    9'd0},{  1'b0, 1'b0, 8'd153,   9'd34},{  1'b0, 1'b0, 8'd152,   9'd80},{  1'b0, 1'b0, 8'd140,    9'd0},{  1'b0, 1'b0, 8'd136,  9'd216},{  1'b0, 1'b0, 8'd121,  9'd348},{  1'b0, 1'b0, 8'd120,    9'd0},{  1'b0, 1'b0, 8'd109,  9'd206},{  1'b0, 1'b0, 8'd109,  9'd214},{  1'b0, 1'b0, 8'd100,    9'd0},{  1'b0, 1'b0,  8'd91,  9'd336},{  1'b0, 1'b0,  8'd83,   9'd22},{  1'b0, 1'b0,  8'd80,    9'd0},{  1'b0, 1'b0,  8'd79,   9'd63},{  1'b0, 1'b0,  8'd77,   9'd30},{  1'b0, 1'b0,  8'd60,    9'd0},{  1'b0, 1'b0,  8'd57,  9'd238},{  1'b0, 1'b0,  8'd50,   9'd37},{  1'b0, 1'b0,  8'd40,    9'd0},{  1'b0, 1'b0,  8'd34,  9'd121},{  1'b0, 1'b0,  8'd25,  9'd312},{  1'b0, 1'b0,  8'd20,    9'd0},{  1'b0, 1'b0,  8'd17,  9'd231},{  1'b0, 1'b0,  8'd15,  9'd196},{  1'b0, 1'b0,   8'd1,  9'd290},{  1'b0, 1'b1,   8'd0,    9'd0},
{  1'b0, 1'b0, 8'd161,    9'd0},{  1'b0, 1'b0, 8'd160,    9'd0},{  1'b0, 1'b0, 8'd156,   9'd84},{  1'b0, 1'b0, 8'd154,   9'd90},{  1'b0, 1'b0, 8'd141,    9'd0},{  1'b0, 1'b0, 8'd137,  9'd198},{  1'b0, 1'b0, 8'd136,  9'd306},{  1'b0, 1'b0, 8'd121,    9'd0},{  1'b0, 1'b0, 8'd115,  9'd330},{  1'b0, 1'b0, 8'd108,  9'd112},{  1'b0, 1'b0, 8'd101,    9'd0},{  1'b0, 1'b0,  8'd92,  9'd226},{  1'b0, 1'b0,  8'd86,   9'd74},{  1'b0, 1'b0,  8'd81,    9'd0},{  1'b0, 1'b0,  8'd66,  9'd291},{  1'b0, 1'b0,  8'd63,   9'd53},{  1'b0, 1'b0,  8'd61,    9'd0},{  1'b0, 1'b0,  8'd59,  9'd307},{  1'b0, 1'b0,  8'd43,   9'd80},{  1'b0, 1'b0,  8'd41,    9'd0},{  1'b0, 1'b0,  8'd35,   9'd49},{  1'b0, 1'b0,  8'd30,  9'd328},{  1'b0, 1'b0,  8'd21,    9'd0},{  1'b0, 1'b0,  8'd17,  9'd119},{  1'b0, 1'b0,   8'd8,  9'd188},{  1'b0, 1'b0,   8'd3,  9'd348},{  1'b0, 1'b1,   8'd1,    9'd0},
{  1'b0, 1'b0, 8'd162,    9'd0},{  1'b0, 1'b0, 8'd161,    9'd0},{  1'b0, 1'b0, 8'd149,  9'd236},{  1'b0, 1'b0, 8'd148,  9'd260},{  1'b0, 1'b0, 8'd142,    9'd0},{  1'b0, 1'b0, 8'd128,  9'd123},{  1'b0, 1'b0, 8'd122,    9'd0},{  1'b0, 1'b0, 8'd122,  9'd353},{  1'b0, 1'b0, 8'd105,  9'd118},{  1'b0, 1'b0, 8'd102,    9'd0},{  1'b0, 1'b0, 8'd101,  9'd103},{  1'b0, 1'b0,  8'd98,   9'd88},{  1'b0, 1'b0,  8'd91,  9'd181},{  1'b0, 1'b0,  8'd82,    9'd0},{  1'b0, 1'b0,  8'd76,  9'd242},{  1'b0, 1'b0,  8'd72,  9'd349},{  1'b0, 1'b0,  8'd62,    9'd0},{  1'b0, 1'b0,  8'd55,  9'd235},{  1'b0, 1'b0,  8'd43,  9'd281},{  1'b0, 1'b0,  8'd42,    9'd0},{  1'b0, 1'b0,  8'd38,  9'd190},{  1'b0, 1'b0,  8'd29,  9'd261},{  1'b0, 1'b0,  8'd22,    9'd0},{  1'b0, 1'b0,  8'd17,   9'd74},{  1'b0, 1'b0,   8'd7,  9'd317},{  1'b0, 1'b0,   8'd2,    9'd0},{  1'b0, 1'b1,   8'd0,  9'd161},
{  1'b0, 1'b0, 8'd163,    9'd0},{  1'b0, 1'b0, 8'd162,    9'd0},{  1'b0, 1'b0, 8'd156,  9'd123},{  1'b0, 1'b0, 8'd145,  9'd202},{  1'b0, 1'b0, 8'd143,    9'd0},{  1'b0, 1'b0, 8'd134,  9'd173},{  1'b0, 1'b0, 8'd131,  9'd312},{  1'b0, 1'b0, 8'd123,    9'd0},{  1'b0, 1'b0, 8'd115,  9'd259},{  1'b0, 1'b0, 8'd114,   9'd70},{  1'b0, 1'b0, 8'd103,    9'd0},{  1'b0, 1'b0,  8'd90,  9'd200},{  1'b0, 1'b0,  8'd83,    9'd0},{  1'b0, 1'b0,  8'd82,   9'd29},{  1'b0, 1'b0,  8'd79,  9'd245},{  1'b0, 1'b0,  8'd63,    9'd0},{  1'b0, 1'b0,  8'd63,  9'd173},{  1'b0, 1'b0,  8'd53,  9'd112},{  1'b0, 1'b0,  8'd45,  9'd289},{  1'b0, 1'b0,  8'd43,    9'd0},{  1'b0, 1'b0,  8'd36,  9'd208},{  1'b0, 1'b0,  8'd26,  9'd117},{  1'b0, 1'b0,  8'd23,    9'd0},{  1'b0, 1'b0,  8'd13,   9'd67},{  1'b0, 1'b0,  8'd13,  9'd296},{  1'b0, 1'b0,   8'd5,  9'd184},{  1'b0, 1'b1,   8'd3,    9'd0},
{  1'b0, 1'b0, 8'd164,    9'd0},{  1'b0, 1'b0, 8'd163,    9'd0},{  1'b0, 1'b0, 8'd158,  9'd214},{  1'b0, 1'b0, 8'd149,  9'd151},{  1'b0, 1'b0, 8'd144,    9'd0},{  1'b0, 1'b0, 8'd132,  9'd132},{  1'b0, 1'b0, 8'd124,    9'd0},{  1'b0, 1'b0, 8'd123,  9'd180},{  1'b0, 1'b0, 8'd119,  9'd338},{  1'b0, 1'b0, 8'd118,  9'd309},{  1'b0, 1'b0, 8'd104,    9'd0},{  1'b0, 1'b0,  8'd93,   9'd58},{  1'b0, 1'b0,  8'd84,    9'd0},{  1'b0, 1'b0,  8'd81,  9'd161},{  1'b0, 1'b0,  8'd74,  9'd248},{  1'b0, 1'b0,  8'd71,  9'd179},{  1'b0, 1'b0,  8'd64,    9'd0},{  1'b0, 1'b0,  8'd51,  9'd147},{  1'b0, 1'b0,  8'd44,    9'd0},{  1'b0, 1'b0,  8'd44,   9'd26},{  1'b0, 1'b0,  8'd24,    9'd0},{  1'b0, 1'b0,  8'd22,   9'd95},{  1'b0, 1'b0,  8'd21,   9'd75},{  1'b0, 1'b0,  8'd16,   9'd82},{  1'b0, 1'b0,   8'd9,   9'd13},{  1'b0, 1'b0,   8'd4,    9'd0},{  1'b0, 1'b1,   8'd4,  9'd313},
{  1'b0, 1'b0, 8'd165,    9'd0},{  1'b0, 1'b0, 8'd164,    9'd0},{  1'b0, 1'b0, 8'd150,  9'd272},{  1'b0, 1'b0, 8'd145,    9'd0},{  1'b0, 1'b0, 8'd144,  9'd194},{  1'b0, 1'b0, 8'd137,   9'd56},{  1'b0, 1'b0, 8'd127,  9'd125},{  1'b0, 1'b0, 8'd125,    9'd0},{  1'b0, 1'b0, 8'd114,   9'd16},{  1'b0, 1'b0, 8'd110,  9'd291},{  1'b0, 1'b0, 8'd105,    9'd0},{  1'b0, 1'b0,  8'd94,   9'd98},{  1'b0, 1'b0,  8'd89,  9'd103},{  1'b0, 1'b0,  8'd85,    9'd0},{  1'b0, 1'b0,  8'd76,  9'd246},{  1'b0, 1'b0,  8'd65,    9'd0},{  1'b0, 1'b0,  8'd61,    9'd7},{  1'b0, 1'b0,  8'd56,  9'd114},{  1'b0, 1'b0,  8'd45,    9'd0},{  1'b0, 1'b0,  8'd44,  9'd300},{  1'b0, 1'b0,  8'd31,  9'd238},{  1'b0, 1'b0,  8'd27,  9'd273},{  1'b0, 1'b0,  8'd25,    9'd0},{  1'b0, 1'b0,  8'd12,  9'd243},{  1'b0, 1'b0,  8'd12,  9'd300},{  1'b0, 1'b0,   8'd5,    9'd0},{  1'b0, 1'b1,   8'd5,  9'd121},
{  1'b0, 1'b0, 8'd166,    9'd0},{  1'b0, 1'b0, 8'd165,    9'd0},{  1'b0, 1'b0, 8'd146,    9'd0},{  1'b0, 1'b0, 8'd144,   9'd72},{  1'b0, 1'b0, 8'd143,  9'd311},{  1'b0, 1'b0, 8'd135,  9'd265},{  1'b0, 1'b0, 8'd128,  9'd240},{  1'b0, 1'b0, 8'd126,    9'd0},{  1'b0, 1'b0, 8'd117,  9'd242},{  1'b0, 1'b0, 8'd106,    9'd0},{  1'b0, 1'b0, 8'd106,   9'd61},{  1'b0, 1'b0,  8'd95,    9'd3},{  1'b0, 1'b0,  8'd86,    9'd0},{  1'b0, 1'b0,  8'd84,  9'd311},{  1'b0, 1'b0,  8'd66,    9'd0},{  1'b0, 1'b0,  8'd61,   9'd65},{  1'b0, 1'b0,  8'd60,  9'd253},{  1'b0, 1'b0,  8'd49,  9'd128},{  1'b0, 1'b0,  8'd46,    9'd0},{  1'b0, 1'b0,  8'd40,  9'd306},{  1'b0, 1'b0,  8'd32,  9'd298},{  1'b0, 1'b0,  8'd26,    9'd0},{  1'b0, 1'b0,  8'd20,  9'd308},{  1'b0, 1'b0,  8'd19,  9'd189},{  1'b0, 1'b0,  8'd12,  9'd164},{  1'b0, 1'b0,   8'd9,  9'd145},{  1'b0, 1'b1,   8'd6,    9'd0},
{  1'b0, 1'b0, 8'd167,    9'd0},{  1'b0, 1'b0, 8'd166,    9'd0},{  1'b0, 1'b0, 8'd147,    9'd0},{  1'b0, 1'b0, 8'd145,  9'd195},{  1'b0, 1'b0, 8'd141,  9'd329},{  1'b0, 1'b0, 8'd131,  9'd331},{  1'b0, 1'b0, 8'd127,    9'd0},{  1'b0, 1'b0, 8'd127,  9'd170},{  1'b0, 1'b0, 8'd119,  9'd356},{  1'b0, 1'b0, 8'd113,  9'd285},{  1'b0, 1'b0, 8'd107,    9'd0},{  1'b0, 1'b0,  8'd88,  9'd105},{  1'b0, 1'b0,  8'd87,    9'd0},{  1'b0, 1'b0,  8'd86,  9'd342},{  1'b0, 1'b0,  8'd70,   9'd50},{  1'b0, 1'b0,  8'd67,    9'd0},{  1'b0, 1'b0,  8'd64,  9'd332},{  1'b0, 1'b0,  8'd59,  9'd176},{  1'b0, 1'b0,  8'd54,   9'd43},{  1'b0, 1'b0,  8'd47,    9'd0},{  1'b0, 1'b0,  8'd27,    9'd0},{  1'b0, 1'b0,  8'd23,  9'd301},{  1'b0, 1'b0,  8'd23,  9'd159},{  1'b0, 1'b0,   8'd9,  9'd296},{  1'b0, 1'b0,   8'd7,    9'd0},{  1'b0, 1'b0,   8'd5,   9'd96},{  1'b0, 1'b1,   8'd2,   9'd46},
{  1'b0, 1'b0, 8'd168,    9'd0},{  1'b0, 1'b0, 8'd167,    9'd0},{  1'b0, 1'b0, 8'd158,  9'd286},{  1'b0, 1'b0, 8'd151,   9'd91},{  1'b0, 1'b0, 8'd148,    9'd0},{  1'b0, 1'b0, 8'd133,  9'd254},{  1'b0, 1'b0, 8'd130,  9'd267},{  1'b0, 1'b0, 8'd128,    9'd0},{  1'b0, 1'b0, 8'd108,    9'd0},{  1'b0, 1'b0, 8'd107,  9'd227},{  1'b0, 1'b0, 8'd103,   9'd61},{  1'b0, 1'b0,  8'd90,  9'd319},{  1'b0, 1'b0,  8'd88,    9'd0},{  1'b0, 1'b0,  8'd82,  9'd151},{  1'b0, 1'b0,  8'd70,  9'd246},{  1'b0, 1'b0,  8'd68,    9'd0},{  1'b0, 1'b0,  8'd60,  9'd107},{  1'b0, 1'b0,  8'd52,  9'd326},{  1'b0, 1'b0,  8'd51,   9'd97},{  1'b0, 1'b0,  8'd48,    9'd0},{  1'b0, 1'b0,  8'd39,  9'd197},{  1'b0, 1'b0,  8'd29,   9'd79},{  1'b0, 1'b0,  8'd28,    9'd0},{  1'b0, 1'b0,   8'd8,    9'd0},{  1'b0, 1'b0,   8'd8,  9'd121},{  1'b0, 1'b0,   8'd1,  9'd267},{  1'b0, 1'b1,   8'd0,  9'd142},
{  1'b0, 1'b0, 8'd169,    9'd0},{  1'b0, 1'b0, 8'd168,    9'd0},{  1'b0, 1'b0, 8'd155,  9'd133},{  1'b0, 1'b0, 8'd149,    9'd0},{  1'b0, 1'b0, 8'd148,  9'd213},{  1'b0, 1'b0, 8'd134,  9'd194},{  1'b0, 1'b0, 8'd129,    9'd0},{  1'b0, 1'b0, 8'd126,  9'd166},{  1'b0, 1'b0, 8'd116,  9'd318},{  1'b0, 1'b0, 8'd116,  9'd228},{  1'b0, 1'b0, 8'd109,    9'd0},{  1'b0, 1'b0,  8'd89,    9'd0},{  1'b0, 1'b0,  8'd88,   9'd82},{  1'b0, 1'b0,  8'd80,  9'd168},{  1'b0, 1'b0,  8'd78,  9'd325},{  1'b0, 1'b0,  8'd72,  9'd143},{  1'b0, 1'b0,  8'd69,    9'd0},{  1'b0, 1'b0,  8'd50,   9'd62},{  1'b0, 1'b0,  8'd49,    9'd0},{  1'b0, 1'b0,  8'd41,   9'd95},{  1'b0, 1'b0,  8'd33,   9'd98},{  1'b0, 1'b0,  8'd33,  9'd193},{  1'b0, 1'b0,  8'd29,    9'd0},{  1'b0, 1'b0,  8'd14,  9'd229},{  1'b0, 1'b0,  8'd13,  9'd176},{  1'b0, 1'b0,   8'd9,    9'd0},{  1'b0, 1'b1,   8'd6,  9'd315},
{  1'b0, 1'b0, 8'd170,    9'd0},{  1'b0, 1'b0, 8'd169,    9'd0},{  1'b0, 1'b0, 8'd154,  9'd334},{  1'b0, 1'b0, 8'd151,   9'd18},{  1'b0, 1'b0, 8'd150,    9'd0},{  1'b0, 1'b0, 8'd130,    9'd0},{  1'b0, 1'b0, 8'd125,    9'd5},{  1'b0, 1'b0, 8'd122,  9'd135},{  1'b0, 1'b0, 8'd110,    9'd0},{  1'b0, 1'b0, 8'd102,  9'd243},{  1'b0, 1'b0, 8'd100,   9'd48},{  1'b0, 1'b0,  8'd96,  9'd148},{  1'b0, 1'b0,  8'd93,  9'd352},{  1'b0, 1'b0,  8'd90,    9'd0},{  1'b0, 1'b0,  8'd75,  9'd220},{  1'b0, 1'b0,  8'd70,    9'd0},{  1'b0, 1'b0,  8'd68,  9'd196},{  1'b0, 1'b0,  8'd50,    9'd0},{  1'b0, 1'b0,  8'd49,  9'd171},{  1'b0, 1'b0,  8'd42,   9'd42},{  1'b0, 1'b0,  8'd30,    9'd0},{  1'b0, 1'b0,  8'd25,  9'd143},{  1'b0, 1'b0,  8'd22,    9'd6},{  1'b0, 1'b0,  8'd10,    9'd0},{  1'b0, 1'b0,  8'd10,   9'd97},{  1'b0, 1'b0,   8'd7,  9'd153},{  1'b0, 1'b1,   8'd2,    9'd4},
{  1'b0, 1'b0, 8'd171,    9'd0},{  1'b0, 1'b0, 8'd170,    9'd0},{  1'b0, 1'b0, 8'd157,  9'd258},{  1'b0, 1'b0, 8'd151,    9'd0},{  1'b0, 1'b0, 8'd142,   9'd55},{  1'b0, 1'b0, 8'd139,  9'd325},{  1'b0, 1'b0, 8'd131,    9'd0},{  1'b0, 1'b0, 8'd120,   9'd97},{  1'b0, 1'b0, 8'd112,  9'd273},{  1'b0, 1'b0, 8'd111,    9'd0},{  1'b0, 1'b0, 8'd107,  9'd345},{  1'b0, 1'b0,  8'd95,  9'd216},{  1'b0, 1'b0,  8'd91,    9'd0},{  1'b0, 1'b0,  8'd80,  9'd151},{  1'b0, 1'b0,  8'd71,    9'd0},{  1'b0, 1'b0,  8'd69,   9'd10},{  1'b0, 1'b0,  8'd62,   9'd43},{  1'b0, 1'b0,  8'd51,    9'd0},{  1'b0, 1'b0,  8'd48,   9'd64},{  1'b0, 1'b0,  8'd45,  9'd262},{  1'b0, 1'b0,  8'd34,  9'd178},{  1'b0, 1'b0,  8'd31,    9'd0},{  1'b0, 1'b0,  8'd26,   9'd65},{  1'b0, 1'b0,  8'd18,  9'd339},{  1'b0, 1'b0,  8'd16,   9'd59},{  1'b0, 1'b0,  8'd11,    9'd0},{  1'b0, 1'b1,  8'd11,  9'd174},
{  1'b0, 1'b0, 8'd172,    9'd0},{  1'b0, 1'b0, 8'd171,    9'd0},{  1'b0, 1'b0, 8'd157,  9'd298},{  1'b0, 1'b0, 8'd152,    9'd0},{  1'b0, 1'b0, 8'd150,  9'd318},{  1'b0, 1'b0, 8'd139,   9'd39},{  1'b0, 1'b0, 8'd133,  9'd210},{  1'b0, 1'b0, 8'd132,    9'd0},{  1'b0, 1'b0, 8'd118,  9'd354},{  1'b0, 1'b0, 8'd112,    9'd0},{  1'b0, 1'b0, 8'd100,  9'd128},{  1'b0, 1'b0,  8'd97,  9'd232},{  1'b0, 1'b0,  8'd92,    9'd0},{  1'b0, 1'b0,  8'd87,   9'd96},{  1'b0, 1'b0,  8'd73,   9'd80},{  1'b0, 1'b0,  8'd72,    9'd0},{  1'b0, 1'b0,  8'd66,  9'd246},{  1'b0, 1'b0,  8'd52,    9'd0},{  1'b0, 1'b0,  8'd46,    9'd8},{  1'b0, 1'b0,  8'd46,  9'd101},{  1'b0, 1'b0,  8'd35,  9'd231},{  1'b0, 1'b0,  8'd32,    9'd0},{  1'b0, 1'b0,  8'd32,  9'd344},{  1'b0, 1'b0,  8'd14,  9'd106},{  1'b0, 1'b0,  8'd12,    9'd0},{  1'b0, 1'b0,   8'd4,   9'd58},{  1'b0, 1'b1,   8'd1,  9'd174},
{  1'b0, 1'b0, 8'd173,    9'd0},{  1'b0, 1'b0, 8'd172,    9'd0},{  1'b0, 1'b0, 8'd153,    9'd0},{  1'b0, 1'b0, 8'd147,   9'd86},{  1'b0, 1'b0, 8'd146,  9'd143},{  1'b0, 1'b0, 8'd133,    9'd0},{  1'b0, 1'b0, 8'd132,  9'd253},{  1'b0, 1'b0, 8'd123,   9'd56},{  1'b0, 1'b0, 8'd113,    9'd0},{  1'b0, 1'b0, 8'd112,  9'd189},{  1'b0, 1'b0, 8'd103,  9'd345},{  1'b0, 1'b0,  8'd94,  9'd180},{  1'b0, 1'b0,  8'd93,    9'd0},{  1'b0, 1'b0,  8'd87,  9'd221},{  1'b0, 1'b0,  8'd74,   9'd47},{  1'b0, 1'b0,  8'd73,    9'd0},{  1'b0, 1'b0,  8'd73,   9'd50},{  1'b0, 1'b0,  8'd54,  9'd186},{  1'b0, 1'b0,  8'd53,    9'd0},{  1'b0, 1'b0,  8'd41,   9'd28},{  1'b0, 1'b0,  8'd37,   9'd48},{  1'b0, 1'b0,  8'd33,    9'd0},{  1'b0, 1'b0,  8'd28,  9'd125},{  1'b0, 1'b0,  8'd13,    9'd0},{  1'b0, 1'b0,  8'd11,  9'd230},{  1'b0, 1'b0,  8'd10,  9'd213},{  1'b0, 1'b1,   8'd8,   9'd30},
{  1'b0, 1'b0, 8'd174,    9'd0},{  1'b0, 1'b0, 8'd173,    9'd0},{  1'b0, 1'b0, 8'd154,    9'd0},{  1'b0, 1'b0, 8'd153,  9'd103},{  1'b0, 1'b0, 8'd140,  9'd196},{  1'b0, 1'b0, 8'd134,    9'd0},{  1'b0, 1'b0, 8'd129,   9'd10},{  1'b0, 1'b0, 8'd124,  9'd184},{  1'b0, 1'b0, 8'd114,    9'd0},{  1'b0, 1'b0, 8'd111,  9'd107},{  1'b0, 1'b0, 8'd110,   9'd23},{  1'b0, 1'b0,  8'd94,    9'd0},{  1'b0, 1'b0,  8'd92,  9'd184},{  1'b0, 1'b0,  8'd85,   9'd54},{  1'b0, 1'b0,  8'd74,    9'd0},{  1'b0, 1'b0,  8'd69,  9'd154},{  1'b0, 1'b0,  8'd64,  9'd277},{  1'b0, 1'b0,  8'd55,   9'd68},{  1'b0, 1'b0,  8'd54,    9'd0},{  1'b0, 1'b0,  8'd42,  9'd201},{  1'b0, 1'b0,  8'd39,  9'd189},{  1'b0, 1'b0,  8'd34,    9'd0},{  1'b0, 1'b0,  8'd31,  9'd102},{  1'b0, 1'b0,  8'd18,  9'd300},{  1'b0, 1'b0,  8'd14,    9'd0},{  1'b0, 1'b0,   8'd7,  9'd357},{  1'b0, 1'b1,   8'd6,  9'd185},
{  1'b0, 1'b0, 8'd175,    9'd0},{  1'b0, 1'b0, 8'd174,    9'd0},{  1'b0, 1'b0, 8'd155,    9'd0},{  1'b0, 1'b0, 8'd152,  9'd234},{  1'b0, 1'b0, 8'd147,  9'd280},{  1'b0, 1'b0, 8'd138,   9'd59},{  1'b0, 1'b0, 8'd135,    9'd0},{  1'b0, 1'b0, 8'd125,   9'd67},{  1'b0, 1'b0, 8'd115,    9'd0},{  1'b0, 1'b0, 8'd113,   9'd79},{  1'b0, 1'b0, 8'd106,   9'd19},{  1'b0, 1'b0,  8'd95,    9'd0},{  1'b0, 1'b0,  8'd85,  9'd244},{  1'b0, 1'b0,  8'd84,  9'd332},{  1'b0, 1'b0,  8'd75,    9'd0},{  1'b0, 1'b0,  8'd75,  9'd227},{  1'b0, 1'b0,  8'd71,   9'd61},{  1'b0, 1'b0,  8'd55,    9'd0},{  1'b0, 1'b0,  8'd47,   9'd93},{  1'b0, 1'b0,  8'd47,  9'd123},{  1'b0, 1'b0,  8'd36,  9'd160},{  1'b0, 1'b0,  8'd35,    9'd0},{  1'b0, 1'b0,  8'd30,   9'd26},{  1'b0, 1'b0,  8'd15,    9'd0},{  1'b0, 1'b0,  8'd14,  9'd201},{  1'b0, 1'b0,   8'd6,  9'd124},{  1'b0, 1'b1,   8'd0,  9'd311},
{  1'b0, 1'b0, 8'd176,    9'd0},{  1'b0, 1'b0, 8'd175,    9'd0},{  1'b0, 1'b0, 8'd159,   9'd84},{  1'b0, 1'b0, 8'd156,    9'd0},{  1'b0, 1'b0, 8'd142,  9'd329},{  1'b0, 1'b0, 8'd136,    9'd0},{  1'b0, 1'b0, 8'd129,  9'd210},{  1'b0, 1'b0, 8'd126,  9'd336},{  1'b0, 1'b0, 8'd117,   9'd44},{  1'b0, 1'b0, 8'd116,    9'd0},{  1'b0, 1'b0, 8'd105,  9'd145},{  1'b0, 1'b0,  8'd99,  9'd286},{  1'b0, 1'b0,  8'd96,    9'd0},{  1'b0, 1'b0,  8'd96,   9'd89},{  1'b0, 1'b0,  8'd76,    9'd0},{  1'b0, 1'b0,  8'd67,  9'd317},{  1'b0, 1'b0,  8'd67,  9'd237},{  1'b0, 1'b0,  8'd56,    9'd0},{  1'b0, 1'b0,  8'd53,  9'd180},{  1'b0, 1'b0,  8'd40,  9'd159},{  1'b0, 1'b0,  8'd36,    9'd0},{  1'b0, 1'b0,  8'd21,  9'd217},{  1'b0, 1'b0,  8'd20,  9'd257},{  1'b0, 1'b0,  8'd18,  9'd329},{  1'b0, 1'b0,  8'd16,    9'd0},{  1'b0, 1'b0,  8'd10,   9'd85},{  1'b0, 1'b1,   8'd3,  9'd225},
{  1'b0, 1'b0, 8'd177,    9'd0},{  1'b0, 1'b0, 8'd176,    9'd0},{  1'b0, 1'b0, 8'd157,    9'd0},{  1'b0, 1'b0, 8'd155,   9'd68},{  1'b0, 1'b0, 8'd143,   9'd72},{  1'b0, 1'b0, 8'd137,    9'd0},{  1'b0, 1'b0, 8'd124,   9'd32},{  1'b0, 1'b0, 8'd121,  9'd155},{  1'b0, 1'b0, 8'd117,    9'd0},{  1'b0, 1'b0, 8'd104,   9'd51},{  1'b0, 1'b0, 8'd102,  9'd229},{  1'b0, 1'b0,  8'd98,  9'd238},{  1'b0, 1'b0,  8'd97,    9'd0},{  1'b0, 1'b0,  8'd81,  9'd177},{  1'b0, 1'b0,  8'd78,  9'd120},{  1'b0, 1'b0,  8'd77,    9'd0},{  1'b0, 1'b0,  8'd65,  9'd291},{  1'b0, 1'b0,  8'd57,    9'd0},{  1'b0, 1'b0,  8'd57,  9'd195},{  1'b0, 1'b0,  8'd48,   9'd24},{  1'b0, 1'b0,  8'd37,    9'd0},{  1'b0, 1'b0,  8'd37,  9'd155},{  1'b0, 1'b0,  8'd28,  9'd330},{  1'b0, 1'b0,  8'd17,    9'd0},{  1'b0, 1'b0,  8'd15,  9'd336},{  1'b0, 1'b0,   8'd4,  9'd161},{  1'b0, 1'b1,   8'd2,  9'd137},
{  1'b0, 1'b0, 8'd178,    9'd0},{  1'b0, 1'b0, 8'd177,    9'd0},{  1'b0, 1'b0, 8'd158,    9'd0},{  1'b0, 1'b0, 8'd141,  9'd161},{  1'b0, 1'b0, 8'd140,  9'd138},{  1'b0, 1'b0, 8'd138,    9'd0},{  1'b0, 1'b0, 8'd135,   9'd23},{  1'b0, 1'b0, 8'd120,  9'd317},{  1'b0, 1'b0, 8'd118,    9'd0},{  1'b0, 1'b0, 8'd111,  9'd277},{  1'b0, 1'b0, 8'd108,  9'd230},{  1'b0, 1'b0,  8'd98,    9'd0},{  1'b0, 1'b0,  8'd97,  9'd160},{  1'b0, 1'b0,  8'd83,  9'd162},{  1'b0, 1'b0,  8'd78,    9'd0},{  1'b0, 1'b0,  8'd77,  9'd288},{  1'b0, 1'b0,  8'd68,   9'd20},{  1'b0, 1'b0,  8'd58,    9'd0},{  1'b0, 1'b0,  8'd58,  9'd202},{  1'b0, 1'b0,  8'd56,  9'd234},{  1'b0, 1'b0,  8'd38,    9'd0},{  1'b0, 1'b0,  8'd38,  9'd309},{  1'b0, 1'b0,  8'd24,  9'd335},{  1'b0, 1'b0,  8'd19,  9'd136},{  1'b0, 1'b0,  8'd19,  9'd295},{  1'b0, 1'b0,  8'd18,    9'd0},{  1'b0, 1'b1,  8'd16,  9'd299},
{  1'b0, 1'b0, 8'd179,    9'd0},{  1'b0, 1'b0, 8'd178,    9'd0},{  1'b0, 1'b0, 8'd159,    9'd0},{  1'b0, 1'b0, 8'd159,   9'd72},{  1'b0, 1'b0, 8'd146,  9'd341},{  1'b0, 1'b0, 8'd139,    9'd0},{  1'b0, 1'b0, 8'd138,  9'd284},{  1'b0, 1'b0, 8'd130,  9'd280},{  1'b0, 1'b0, 8'd119,    9'd0},{  1'b0, 1'b0, 8'd104,  9'd207},{  1'b0, 1'b0, 8'd101,  9'd329},{  1'b0, 1'b0,  8'd99,    9'd0},{  1'b0, 1'b0,  8'd99,   9'd69},{  1'b0, 1'b0,  8'd89,  9'd105},{  1'b0, 1'b0,  8'd79,    9'd0},{  1'b0, 1'b0,  8'd65,   9'd16},{  1'b0, 1'b0,  8'd62,  9'd115},{  1'b0, 1'b0,  8'd59,    9'd0},{  1'b0, 1'b0,  8'd58,   9'd92},{  1'b0, 1'b0,  8'd52,  9'd144},{  1'b0, 1'b0,  8'd39,    9'd0},{  1'b0, 1'b0,  8'd27,   9'd51},{  1'b0, 1'b0,  8'd24,   9'd37},{  1'b0, 1'b0,  8'd19,    9'd0},{  1'b0, 1'b0,  8'd15,   9'd78},{  1'b0, 1'b0,  8'd11,  9'd308},{  1'b0, 1'b1,   8'd3,  9'd236}
};
localparam bit [18 : 0] cLARGE_HS_V_TAB_8BY9_PACKED[cLARGE_HS_TAB_8BY9_PACKED_SIZE] = '{
{8'd179, 1'b0,   10'd0},{8'd179, 1'b1, 10'd513},
{8'd178, 1'b0, 10'd486},{8'd178, 1'b1, 10'd514},
{8'd177, 1'b0, 10'd459},{8'd177, 1'b1, 10'd487},
{8'd176, 1'b0, 10'd432},{8'd176, 1'b1, 10'd460},
{8'd175, 1'b0, 10'd405},{8'd175, 1'b1, 10'd433},
{8'd174, 1'b0, 10'd378},{8'd174, 1'b1, 10'd406},
{8'd173, 1'b0, 10'd351},{8'd173, 1'b1, 10'd379},
{8'd172, 1'b0, 10'd324},{8'd172, 1'b1, 10'd352},
{8'd171, 1'b0, 10'd297},{8'd171, 1'b1, 10'd325},
{8'd170, 1'b0, 10'd270},{8'd170, 1'b1, 10'd298},
{8'd169, 1'b0, 10'd243},{8'd169, 1'b1, 10'd271},
{8'd168, 1'b0, 10'd216},{8'd168, 1'b1, 10'd244},
{8'd167, 1'b0, 10'd189},{8'd167, 1'b1, 10'd217},
{8'd166, 1'b0, 10'd162},{8'd166, 1'b1, 10'd190},
{8'd165, 1'b0, 10'd135},{8'd165, 1'b1, 10'd163},
{8'd164, 1'b0, 10'd108},{8'd164, 1'b1, 10'd136},
{8'd163, 1'b0,  10'd81},{8'd163, 1'b1, 10'd109},
{8'd162, 1'b0,  10'd54},{8'd162, 1'b1,  10'd82},
{8'd161, 1'b0,  10'd27},{8'd161, 1'b1,  10'd55},
{8'd160, 1'b0,   10'd1},{8'd160, 1'b1,  10'd28},
{8'd159, 1'b0, 10'd434},{8'd159, 1'b0, 10'd515},{8'd159, 1'b1, 10'd516},
{8'd158, 1'b0, 10'd110},{8'd158, 1'b0, 10'd218},{8'd158, 1'b1, 10'd488},
{8'd157, 1'b0, 10'd299},{8'd157, 1'b0, 10'd326},{8'd157, 1'b1, 10'd461},
{8'd156, 1'b0,  10'd29},{8'd156, 1'b0,  10'd83},{8'd156, 1'b1, 10'd435},
{8'd155, 1'b0, 10'd245},{8'd155, 1'b0, 10'd407},{8'd155, 1'b1, 10'd462},
{8'd154, 1'b0,  10'd30},{8'd154, 1'b0, 10'd272},{8'd154, 1'b1, 10'd380},
{8'd153, 1'b0,   10'd2},{8'd153, 1'b0, 10'd353},{8'd153, 1'b1, 10'd381},
{8'd152, 1'b0,   10'd3},{8'd152, 1'b0, 10'd327},{8'd152, 1'b1, 10'd408},
{8'd151, 1'b0, 10'd219},{8'd151, 1'b0, 10'd273},{8'd151, 1'b1, 10'd300},
{8'd150, 1'b0, 10'd137},{8'd150, 1'b0, 10'd274},{8'd150, 1'b1, 10'd328},
{8'd149, 1'b0,  10'd56},{8'd149, 1'b0, 10'd111},{8'd149, 1'b1, 10'd246},
{8'd148, 1'b0,  10'd57},{8'd148, 1'b0, 10'd220},{8'd148, 1'b1, 10'd247},
{8'd147, 1'b0, 10'd191},{8'd147, 1'b0, 10'd354},{8'd147, 1'b1, 10'd409},
{8'd146, 1'b0, 10'd164},{8'd146, 1'b0, 10'd355},{8'd146, 1'b1, 10'd517},
{8'd145, 1'b0,  10'd84},{8'd145, 1'b0, 10'd138},{8'd145, 1'b1, 10'd192},
{8'd144, 1'b0, 10'd112},{8'd144, 1'b0, 10'd139},{8'd144, 1'b1, 10'd165},
{8'd143, 1'b0,  10'd85},{8'd143, 1'b0, 10'd166},{8'd143, 1'b1, 10'd463},
{8'd142, 1'b0,  10'd58},{8'd142, 1'b0, 10'd301},{8'd142, 1'b1, 10'd436},
{8'd141, 1'b0,  10'd31},{8'd141, 1'b0, 10'd193},{8'd141, 1'b1, 10'd489},
{8'd140, 1'b0,   10'd4},{8'd140, 1'b0, 10'd382},{8'd140, 1'b1, 10'd490},
{8'd139, 1'b0, 10'd302},{8'd139, 1'b0, 10'd329},{8'd139, 1'b1, 10'd518},
{8'd138, 1'b0, 10'd410},{8'd138, 1'b0, 10'd491},{8'd138, 1'b1, 10'd519},
{8'd137, 1'b0,  10'd32},{8'd137, 1'b0, 10'd140},{8'd137, 1'b1, 10'd464},
{8'd136, 1'b0,   10'd5},{8'd136, 1'b0,  10'd33},{8'd136, 1'b1, 10'd437},
{8'd135, 1'b0, 10'd167},{8'd135, 1'b0, 10'd411},{8'd135, 1'b1, 10'd492},
{8'd134, 1'b0,  10'd86},{8'd134, 1'b0, 10'd248},{8'd134, 1'b1, 10'd383},
{8'd133, 1'b0, 10'd221},{8'd133, 1'b0, 10'd330},{8'd133, 1'b1, 10'd356},
{8'd132, 1'b0, 10'd113},{8'd132, 1'b0, 10'd331},{8'd132, 1'b1, 10'd357},
{8'd131, 1'b0,  10'd87},{8'd131, 1'b0, 10'd194},{8'd131, 1'b1, 10'd303},
{8'd130, 1'b0, 10'd222},{8'd130, 1'b0, 10'd275},{8'd130, 1'b1, 10'd520},
{8'd129, 1'b0, 10'd249},{8'd129, 1'b0, 10'd384},{8'd129, 1'b1, 10'd438},
{8'd128, 1'b0,  10'd59},{8'd128, 1'b0, 10'd168},{8'd128, 1'b1, 10'd223},
{8'd127, 1'b0, 10'd141},{8'd127, 1'b0, 10'd195},{8'd127, 1'b1, 10'd196},
{8'd126, 1'b0, 10'd169},{8'd126, 1'b0, 10'd250},{8'd126, 1'b1, 10'd439},
{8'd125, 1'b0, 10'd142},{8'd125, 1'b0, 10'd276},{8'd125, 1'b1, 10'd412},
{8'd124, 1'b0, 10'd114},{8'd124, 1'b0, 10'd385},{8'd124, 1'b1, 10'd465},
{8'd123, 1'b0,  10'd88},{8'd123, 1'b0, 10'd115},{8'd123, 1'b1, 10'd358},
{8'd122, 1'b0,  10'd60},{8'd122, 1'b0,  10'd61},{8'd122, 1'b1, 10'd277},
{8'd121, 1'b0,   10'd6},{8'd121, 1'b0,  10'd34},{8'd121, 1'b1, 10'd466},
{8'd120, 1'b0,   10'd7},{8'd120, 1'b0, 10'd304},{8'd120, 1'b1, 10'd493},
{8'd119, 1'b0, 10'd116},{8'd119, 1'b0, 10'd197},{8'd119, 1'b1, 10'd521},
{8'd118, 1'b0, 10'd117},{8'd118, 1'b0, 10'd332},{8'd118, 1'b1, 10'd494},
{8'd117, 1'b0, 10'd170},{8'd117, 1'b0, 10'd440},{8'd117, 1'b1, 10'd467},
{8'd116, 1'b0, 10'd251},{8'd116, 1'b0, 10'd252},{8'd116, 1'b1, 10'd441},
{8'd115, 1'b0,  10'd35},{8'd115, 1'b0,  10'd89},{8'd115, 1'b1, 10'd413},
{8'd114, 1'b0,  10'd90},{8'd114, 1'b0, 10'd143},{8'd114, 1'b1, 10'd386},
{8'd113, 1'b0, 10'd198},{8'd113, 1'b0, 10'd359},{8'd113, 1'b1, 10'd414},
{8'd112, 1'b0, 10'd305},{8'd112, 1'b0, 10'd333},{8'd112, 1'b1, 10'd360},
{8'd111, 1'b0, 10'd306},{8'd111, 1'b0, 10'd387},{8'd111, 1'b1, 10'd495},
{8'd110, 1'b0, 10'd144},{8'd110, 1'b0, 10'd278},{8'd110, 1'b1, 10'd388},
{8'd109, 1'b0,   10'd8},{8'd109, 1'b0,   10'd9},{8'd109, 1'b1, 10'd253},
{8'd108, 1'b0,  10'd36},{8'd108, 1'b0, 10'd224},{8'd108, 1'b1, 10'd496},
{8'd107, 1'b0, 10'd199},{8'd107, 1'b0, 10'd225},{8'd107, 1'b1, 10'd307},
{8'd106, 1'b0, 10'd171},{8'd106, 1'b0, 10'd172},{8'd106, 1'b1, 10'd415},
{8'd105, 1'b0,  10'd62},{8'd105, 1'b0, 10'd145},{8'd105, 1'b1, 10'd442},
{8'd104, 1'b0, 10'd118},{8'd104, 1'b0, 10'd468},{8'd104, 1'b1, 10'd522},
{8'd103, 1'b0,  10'd91},{8'd103, 1'b0, 10'd226},{8'd103, 1'b1, 10'd361},
{8'd102, 1'b0,  10'd63},{8'd102, 1'b0, 10'd279},{8'd102, 1'b1, 10'd469},
{8'd101, 1'b0,  10'd37},{8'd101, 1'b0,  10'd64},{8'd101, 1'b1, 10'd523},
{8'd100, 1'b0,  10'd10},{8'd100, 1'b0, 10'd280},{8'd100, 1'b1, 10'd334},
{ 8'd99, 1'b0, 10'd443},{ 8'd99, 1'b0, 10'd524},{ 8'd99, 1'b1, 10'd525},
{ 8'd98, 1'b0,  10'd65},{ 8'd98, 1'b0, 10'd470},{ 8'd98, 1'b1, 10'd497},
{ 8'd97, 1'b0, 10'd335},{ 8'd97, 1'b0, 10'd471},{ 8'd97, 1'b1, 10'd498},
{ 8'd96, 1'b0, 10'd281},{ 8'd96, 1'b0, 10'd444},{ 8'd96, 1'b1, 10'd445},
{ 8'd95, 1'b0, 10'd173},{ 8'd95, 1'b0, 10'd308},{ 8'd95, 1'b1, 10'd416},
{ 8'd94, 1'b0, 10'd146},{ 8'd94, 1'b0, 10'd362},{ 8'd94, 1'b1, 10'd389},
{ 8'd93, 1'b0, 10'd119},{ 8'd93, 1'b0, 10'd282},{ 8'd93, 1'b1, 10'd363},
{ 8'd92, 1'b0,  10'd38},{ 8'd92, 1'b0, 10'd336},{ 8'd92, 1'b1, 10'd390},
{ 8'd91, 1'b0,  10'd11},{ 8'd91, 1'b0,  10'd66},{ 8'd91, 1'b1, 10'd309},
{ 8'd90, 1'b0,  10'd92},{ 8'd90, 1'b0, 10'd227},{ 8'd90, 1'b1, 10'd283},
{ 8'd89, 1'b0, 10'd147},{ 8'd89, 1'b0, 10'd254},{ 8'd89, 1'b1, 10'd526},
{ 8'd88, 1'b0, 10'd200},{ 8'd88, 1'b0, 10'd228},{ 8'd88, 1'b1, 10'd255},
{ 8'd87, 1'b0, 10'd201},{ 8'd87, 1'b0, 10'd337},{ 8'd87, 1'b1, 10'd364},
{ 8'd86, 1'b0,  10'd39},{ 8'd86, 1'b0, 10'd174},{ 8'd86, 1'b1, 10'd202},
{ 8'd85, 1'b0, 10'd148},{ 8'd85, 1'b0, 10'd391},{ 8'd85, 1'b1, 10'd417},
{ 8'd84, 1'b0, 10'd120},{ 8'd84, 1'b0, 10'd175},{ 8'd84, 1'b1, 10'd418},
{ 8'd83, 1'b0,  10'd12},{ 8'd83, 1'b0,  10'd93},{ 8'd83, 1'b1, 10'd499},
{ 8'd82, 1'b0,  10'd67},{ 8'd82, 1'b0,  10'd94},{ 8'd82, 1'b1, 10'd229},
{ 8'd81, 1'b0,  10'd40},{ 8'd81, 1'b0, 10'd121},{ 8'd81, 1'b1, 10'd472},
{ 8'd80, 1'b0,  10'd13},{ 8'd80, 1'b0, 10'd256},{ 8'd80, 1'b1, 10'd310},
{ 8'd79, 1'b0,  10'd14},{ 8'd79, 1'b0,  10'd95},{ 8'd79, 1'b1, 10'd527},
{ 8'd78, 1'b0, 10'd257},{ 8'd78, 1'b0, 10'd473},{ 8'd78, 1'b1, 10'd500},
{ 8'd77, 1'b0,  10'd15},{ 8'd77, 1'b0, 10'd474},{ 8'd77, 1'b1, 10'd501},
{ 8'd76, 1'b0,  10'd68},{ 8'd76, 1'b0, 10'd149},{ 8'd76, 1'b1, 10'd446},
{ 8'd75, 1'b0, 10'd284},{ 8'd75, 1'b0, 10'd419},{ 8'd75, 1'b1, 10'd420},
{ 8'd74, 1'b0, 10'd122},{ 8'd74, 1'b0, 10'd365},{ 8'd74, 1'b1, 10'd392},
{ 8'd73, 1'b0, 10'd338},{ 8'd73, 1'b0, 10'd366},{ 8'd73, 1'b1, 10'd367},
{ 8'd72, 1'b0,  10'd69},{ 8'd72, 1'b0, 10'd258},{ 8'd72, 1'b1, 10'd339},
{ 8'd71, 1'b0, 10'd123},{ 8'd71, 1'b0, 10'd311},{ 8'd71, 1'b1, 10'd421},
{ 8'd70, 1'b0, 10'd203},{ 8'd70, 1'b0, 10'd230},{ 8'd70, 1'b1, 10'd285},
{ 8'd69, 1'b0, 10'd259},{ 8'd69, 1'b0, 10'd312},{ 8'd69, 1'b1, 10'd393},
{ 8'd68, 1'b0, 10'd231},{ 8'd68, 1'b0, 10'd286},{ 8'd68, 1'b1, 10'd502},
{ 8'd67, 1'b0, 10'd204},{ 8'd67, 1'b0, 10'd447},{ 8'd67, 1'b1, 10'd448},
{ 8'd66, 1'b0,  10'd41},{ 8'd66, 1'b0, 10'd176},{ 8'd66, 1'b1, 10'd340},
{ 8'd65, 1'b0, 10'd150},{ 8'd65, 1'b0, 10'd475},{ 8'd65, 1'b1, 10'd528},
{ 8'd64, 1'b0, 10'd124},{ 8'd64, 1'b0, 10'd205},{ 8'd64, 1'b1, 10'd394},
{ 8'd63, 1'b0,  10'd42},{ 8'd63, 1'b0,  10'd96},{ 8'd63, 1'b1,  10'd97},
{ 8'd62, 1'b0,  10'd70},{ 8'd62, 1'b0, 10'd313},{ 8'd62, 1'b1, 10'd529},
{ 8'd61, 1'b0,  10'd43},{ 8'd61, 1'b0, 10'd151},{ 8'd61, 1'b1, 10'd177},
{ 8'd60, 1'b0,  10'd16},{ 8'd60, 1'b0, 10'd178},{ 8'd60, 1'b1, 10'd232},
{ 8'd59, 1'b0,  10'd44},{ 8'd59, 1'b0, 10'd206},{ 8'd59, 1'b1, 10'd530},
{ 8'd58, 1'b0, 10'd503},{ 8'd58, 1'b0, 10'd504},{ 8'd58, 1'b1, 10'd531},
{ 8'd57, 1'b0,  10'd17},{ 8'd57, 1'b0, 10'd476},{ 8'd57, 1'b1, 10'd477},
{ 8'd56, 1'b0, 10'd152},{ 8'd56, 1'b0, 10'd449},{ 8'd56, 1'b1, 10'd505},
{ 8'd55, 1'b0,  10'd71},{ 8'd55, 1'b0, 10'd395},{ 8'd55, 1'b1, 10'd422},
{ 8'd54, 1'b0, 10'd207},{ 8'd54, 1'b0, 10'd368},{ 8'd54, 1'b1, 10'd396},
{ 8'd53, 1'b0,  10'd98},{ 8'd53, 1'b0, 10'd369},{ 8'd53, 1'b1, 10'd450},
{ 8'd52, 1'b0, 10'd233},{ 8'd52, 1'b0, 10'd341},{ 8'd52, 1'b1, 10'd532},
{ 8'd51, 1'b0, 10'd125},{ 8'd51, 1'b0, 10'd234},{ 8'd51, 1'b1, 10'd314},
{ 8'd50, 1'b0,  10'd18},{ 8'd50, 1'b0, 10'd260},{ 8'd50, 1'b1, 10'd287},
{ 8'd49, 1'b0, 10'd179},{ 8'd49, 1'b0, 10'd261},{ 8'd49, 1'b1, 10'd288},
{ 8'd48, 1'b0, 10'd235},{ 8'd48, 1'b0, 10'd315},{ 8'd48, 1'b1, 10'd478},
{ 8'd47, 1'b0, 10'd208},{ 8'd47, 1'b0, 10'd423},{ 8'd47, 1'b1, 10'd424},
{ 8'd46, 1'b0, 10'd180},{ 8'd46, 1'b0, 10'd342},{ 8'd46, 1'b1, 10'd343},
{ 8'd45, 1'b0,  10'd99},{ 8'd45, 1'b0, 10'd153},{ 8'd45, 1'b1, 10'd316},
{ 8'd44, 1'b0, 10'd126},{ 8'd44, 1'b0, 10'd127},{ 8'd44, 1'b1, 10'd154},
{ 8'd43, 1'b0,  10'd45},{ 8'd43, 1'b0,  10'd72},{ 8'd43, 1'b1, 10'd100},
{ 8'd42, 1'b0,  10'd73},{ 8'd42, 1'b0, 10'd289},{ 8'd42, 1'b1, 10'd397},
{ 8'd41, 1'b0,  10'd46},{ 8'd41, 1'b0, 10'd262},{ 8'd41, 1'b1, 10'd370},
{ 8'd40, 1'b0,  10'd19},{ 8'd40, 1'b0, 10'd181},{ 8'd40, 1'b1, 10'd451},
{ 8'd39, 1'b0, 10'd236},{ 8'd39, 1'b0, 10'd398},{ 8'd39, 1'b1, 10'd533},
{ 8'd38, 1'b0,  10'd74},{ 8'd38, 1'b0, 10'd506},{ 8'd38, 1'b1, 10'd507},
{ 8'd37, 1'b0, 10'd371},{ 8'd37, 1'b0, 10'd479},{ 8'd37, 1'b1, 10'd480},
{ 8'd36, 1'b0, 10'd101},{ 8'd36, 1'b0, 10'd425},{ 8'd36, 1'b1, 10'd452},
{ 8'd35, 1'b0,  10'd47},{ 8'd35, 1'b0, 10'd344},{ 8'd35, 1'b1, 10'd426},
{ 8'd34, 1'b0,  10'd20},{ 8'd34, 1'b0, 10'd317},{ 8'd34, 1'b1, 10'd399},
{ 8'd33, 1'b0, 10'd263},{ 8'd33, 1'b0, 10'd264},{ 8'd33, 1'b1, 10'd372},
{ 8'd32, 1'b0, 10'd182},{ 8'd32, 1'b0, 10'd345},{ 8'd32, 1'b1, 10'd346},
{ 8'd31, 1'b0, 10'd155},{ 8'd31, 1'b0, 10'd318},{ 8'd31, 1'b1, 10'd400},
{ 8'd30, 1'b0,  10'd48},{ 8'd30, 1'b0, 10'd290},{ 8'd30, 1'b1, 10'd427},
{ 8'd29, 1'b0,  10'd75},{ 8'd29, 1'b0, 10'd237},{ 8'd29, 1'b1, 10'd265},
{ 8'd28, 1'b0, 10'd238},{ 8'd28, 1'b0, 10'd373},{ 8'd28, 1'b1, 10'd481},
{ 8'd27, 1'b0, 10'd156},{ 8'd27, 1'b0, 10'd209},{ 8'd27, 1'b1, 10'd534},
{ 8'd26, 1'b0, 10'd102},{ 8'd26, 1'b0, 10'd183},{ 8'd26, 1'b1, 10'd319},
{ 8'd25, 1'b0,  10'd21},{ 8'd25, 1'b0, 10'd157},{ 8'd25, 1'b1, 10'd291},
{ 8'd24, 1'b0, 10'd128},{ 8'd24, 1'b0, 10'd508},{ 8'd24, 1'b1, 10'd535},
{ 8'd23, 1'b0, 10'd103},{ 8'd23, 1'b0, 10'd210},{ 8'd23, 1'b1, 10'd211},
{ 8'd22, 1'b0,  10'd76},{ 8'd22, 1'b0, 10'd129},{ 8'd22, 1'b1, 10'd292},
{ 8'd21, 1'b0,  10'd49},{ 8'd21, 1'b0, 10'd130},{ 8'd21, 1'b1, 10'd453},
{ 8'd20, 1'b0,  10'd22},{ 8'd20, 1'b0, 10'd184},{ 8'd20, 1'b1, 10'd454},
{ 8'd19, 1'b0, 10'd185},{ 8'd19, 1'b0, 10'd509},{ 8'd19, 1'b0, 10'd510},{ 8'd19, 1'b1, 10'd536},
{ 8'd18, 1'b0, 10'd320},{ 8'd18, 1'b0, 10'd401},{ 8'd18, 1'b0, 10'd455},{ 8'd18, 1'b1, 10'd511},
{ 8'd17, 1'b0,  10'd23},{ 8'd17, 1'b0,  10'd50},{ 8'd17, 1'b0,  10'd77},{ 8'd17, 1'b1, 10'd482},
{ 8'd16, 1'b0, 10'd131},{ 8'd16, 1'b0, 10'd321},{ 8'd16, 1'b0, 10'd456},{ 8'd16, 1'b1, 10'd512},
{ 8'd15, 1'b0,  10'd24},{ 8'd15, 1'b0, 10'd428},{ 8'd15, 1'b0, 10'd483},{ 8'd15, 1'b1, 10'd537},
{ 8'd14, 1'b0, 10'd266},{ 8'd14, 1'b0, 10'd347},{ 8'd14, 1'b0, 10'd402},{ 8'd14, 1'b1, 10'd429},
{ 8'd13, 1'b0, 10'd104},{ 8'd13, 1'b0, 10'd105},{ 8'd13, 1'b0, 10'd267},{ 8'd13, 1'b1, 10'd374},
{ 8'd12, 1'b0, 10'd158},{ 8'd12, 1'b0, 10'd159},{ 8'd12, 1'b0, 10'd186},{ 8'd12, 1'b1, 10'd348},
{ 8'd11, 1'b0, 10'd322},{ 8'd11, 1'b0, 10'd323},{ 8'd11, 1'b0, 10'd375},{ 8'd11, 1'b1, 10'd538},
{ 8'd10, 1'b0, 10'd293},{ 8'd10, 1'b0, 10'd294},{ 8'd10, 1'b0, 10'd376},{ 8'd10, 1'b1, 10'd457},
{  8'd9, 1'b0, 10'd132},{  8'd9, 1'b0, 10'd187},{  8'd9, 1'b0, 10'd212},{  8'd9, 1'b1, 10'd268},
{  8'd8, 1'b0,  10'd51},{  8'd8, 1'b0, 10'd239},{  8'd8, 1'b0, 10'd240},{  8'd8, 1'b1, 10'd377},
{  8'd7, 1'b0,  10'd78},{  8'd7, 1'b0, 10'd213},{  8'd7, 1'b0, 10'd295},{  8'd7, 1'b1, 10'd403},
{  8'd6, 1'b0, 10'd188},{  8'd6, 1'b0, 10'd269},{  8'd6, 1'b0, 10'd404},{  8'd6, 1'b1, 10'd430},
{  8'd5, 1'b0, 10'd106},{  8'd5, 1'b0, 10'd160},{  8'd5, 1'b0, 10'd161},{  8'd5, 1'b1, 10'd214},
{  8'd4, 1'b0, 10'd133},{  8'd4, 1'b0, 10'd134},{  8'd4, 1'b0, 10'd349},{  8'd4, 1'b1, 10'd484},
{  8'd3, 1'b0,  10'd52},{  8'd3, 1'b0, 10'd107},{  8'd3, 1'b0, 10'd458},{  8'd3, 1'b1, 10'd539},
{  8'd2, 1'b0,  10'd79},{  8'd2, 1'b0, 10'd215},{  8'd2, 1'b0, 10'd296},{  8'd2, 1'b1, 10'd485},
{  8'd1, 1'b0,  10'd25},{  8'd1, 1'b0,  10'd53},{  8'd1, 1'b0, 10'd241},{  8'd1, 1'b1, 10'd350},
{  8'd0, 1'b0,  10'd26},{  8'd0, 1'b0,  10'd80},{  8'd0, 1'b0, 10'd242},{  8'd0, 1'b1, 10'd431}
};
localparam int          cLARGE_HS_TAB_9BY10_PACKED_SIZE = 540;
localparam bit [18 : 0] cLARGE_HS_TAB_9BY10_PACKED[cLARGE_HS_TAB_9BY10_PACKED_SIZE] = '{
{  1'b1, 1'b0, 8'd179,    9'd1},{  1'b0, 1'b0, 8'd162,    9'd0},{  1'b0, 1'b0, 8'd154,   9'd64},{  1'b0, 1'b0, 8'd153,   9'd65},{  1'b0, 1'b0, 8'd144,    9'd0},{  1'b0, 1'b0, 8'd131,   9'd58},{  1'b0, 1'b0, 8'd126,    9'd0},{  1'b0, 1'b0, 8'd126,   9'd94},{  1'b0, 1'b0, 8'd124,  9'd216},{  1'b0, 1'b0, 8'd112,  9'd348},{  1'b0, 1'b0, 8'd108,    9'd0},{  1'b0, 1'b0,  8'd97,  9'd237},{  1'b0, 1'b0,  8'd91,    9'd8},{  1'b0, 1'b0,  8'd90,    9'd0},{  1'b0, 1'b0,  8'd86,  9'd103},{  1'b0, 1'b0,  8'd84,   9'd74},{  1'b0, 1'b0,  8'd72,    9'd0},{  1'b0, 1'b0,  8'd64,  9'd291},{  1'b0, 1'b0,  8'd57,  9'd114},{  1'b0, 1'b0,  8'd54,    9'd0},{  1'b0, 1'b0,  8'd53,  9'd126},{  1'b0, 1'b0,  8'd37,  9'd208},{  1'b0, 1'b0,  8'd36,    9'd0},{  1'b0, 1'b0,  8'd35,  9'd121},{  1'b0, 1'b0,  8'd26,  9'd312},{  1'b0, 1'b0,  8'd18,    9'd0},{  1'b0, 1'b0,  8'd13,  9'd196},{  1'b0, 1'b0,  8'd11,  9'd300},{  1'b0, 1'b0,   8'd1,  9'd290},{  1'b0, 1'b1,   8'd0,    9'd0},
{  1'b0, 1'b0, 8'd163,    9'd0},{  1'b0, 1'b0, 8'd162,    9'd0},{  1'b0, 1'b0, 8'd158,  9'd300},{  1'b0, 1'b0, 8'd145,    9'd0},{  1'b0, 1'b0, 8'd144,  9'd321},{  1'b0, 1'b0, 8'd143,  9'd234},{  1'b0, 1'b0, 8'd140,   9'd36},{  1'b0, 1'b0, 8'd127,    9'd0},{  1'b0, 1'b0, 8'd119,   9'd36},{  1'b0, 1'b0, 8'd118,  9'd296},{  1'b0, 1'b0, 8'd109,    9'd0},{  1'b0, 1'b0, 8'd100,  9'd214},{  1'b0, 1'b0,  8'd94,  9'd103},{  1'b0, 1'b0,  8'd91,    9'd0},{  1'b0, 1'b0,  8'd87,  9'd200},{  1'b0, 1'b0,  8'd75,   9'd30},{  1'b0, 1'b0,  8'd73,    9'd0},{  1'b0, 1'b0,  8'd62,  9'd173},{  1'b0, 1'b0,  8'd56,  9'd235},{  1'b0, 1'b0,  8'd55,    9'd0},{  1'b0, 1'b0,  8'd44,  9'd281},{  1'b0, 1'b0,  8'd44,   9'd80},{  1'b0, 1'b0,  8'd37,    9'd0},{  1'b0, 1'b0,  8'd31,  9'd328},{  1'b0, 1'b0,  8'd30,  9'd261},{  1'b0, 1'b0,  8'd19,    9'd0},{  1'b0, 1'b0,  8'd12,  9'd296},{  1'b0, 1'b0,   8'd7,  9'd188},{  1'b0, 1'b0,   8'd3,  9'd348},{  1'b0, 1'b1,   8'd1,    9'd0},
{  1'b0, 1'b0, 8'd164,    9'd0},{  1'b0, 1'b0, 8'd163,    9'd0},{  1'b0, 1'b0, 8'd159,  9'd282},{  1'b0, 1'b0, 8'd146,    9'd0},{  1'b0, 1'b0, 8'd146,   9'd84},{  1'b0, 1'b0, 8'd143,   9'd80},{  1'b0, 1'b0, 8'd137,  9'd260},{  1'b0, 1'b0, 8'd128,    9'd0},{  1'b0, 1'b0, 8'd124,  9'd306},{  1'b0, 1'b0, 8'd110,    9'd0},{  1'b0, 1'b0, 8'd109,  9'd289},{  1'b0, 1'b0, 8'd100,  9'd206},{  1'b0, 1'b0,  8'd98,  9'd112},{  1'b0, 1'b0,  8'd92,    9'd0},{  1'b0, 1'b0,  8'd82,  9'd243},{  1'b0, 1'b0,  8'd79,  9'd229},{  1'b0, 1'b0,  8'd74,    9'd0},{  1'b0, 1'b0,  8'd62,   9'd53},{  1'b0, 1'b0,  8'd58,  9'd238},{  1'b0, 1'b0,  8'd56,    9'd0},{  1'b0, 1'b0,  8'd40,  9'd189},{  1'b0, 1'b0,  8'd38,    9'd0},{  1'b0, 1'b0,  8'd36,   9'd49},{  1'b0, 1'b0,  8'd34,  9'd193},{  1'b0, 1'b0,  8'd27,  9'd117},{  1'b0, 1'b0,  8'd20,    9'd0},{  1'b0, 1'b0,  8'd16,   9'd74},{  1'b0, 1'b0,   8'd8,   9'd13},{  1'b0, 1'b0,   8'd2,    9'd0},{  1'b0, 1'b1,   8'd0,  9'd161},
{  1'b0, 1'b0, 8'd165,    9'd0},{  1'b0, 1'b0, 8'd164,    9'd0},{  1'b0, 1'b0, 8'd152,   9'd75},{  1'b0, 1'b0, 8'd147,    9'd0},{  1'b0, 1'b0, 8'd146,  9'd123},{  1'b0, 1'b0, 8'd138,  9'd169},{  1'b0, 1'b0, 8'd135,  9'd202},{  1'b0, 1'b0, 8'd129,    9'd0},{  1'b0, 1'b0, 8'd111,    9'd0},{  1'b0, 1'b0, 8'd110,  9'd309},{  1'b0, 1'b0, 8'd108,  9'd176},{  1'b0, 1'b0, 8'd106,  9'd259},{  1'b0, 1'b0, 8'd105,   9'd70},{  1'b0, 1'b0,  8'd93,    9'd0},{  1'b0, 1'b0,  8'd79,   9'd60},{  1'b0, 1'b0,  8'd78,   9'd29},{  1'b0, 1'b0,  8'd75,    9'd0},{  1'b0, 1'b0,  8'd71,   9'd50},{  1'b0, 1'b0,  8'd69,  9'd179},{  1'b0, 1'b0,  8'd57,    9'd0},{  1'b0, 1'b0,  8'd52,   9'd37},{  1'b0, 1'b0,  8'd39,    9'd0},{  1'b0, 1'b0,  8'd39,  9'd190},{  1'b0, 1'b0,  8'd23,   9'd95},{  1'b0, 1'b0,  8'd21,    9'd0},{  1'b0, 1'b0,  8'd20,  9'd189},{  1'b0, 1'b0,  8'd16,  9'd119},{  1'b0, 1'b0,  8'd12,   9'd67},{  1'b0, 1'b0,   8'd5,  9'd184},{  1'b0, 1'b1,   8'd3,    9'd0},
{  1'b0, 1'b0, 8'd166,    9'd0},{  1'b0, 1'b0, 8'd165,    9'd0},{  1'b0, 1'b0, 8'd155,  9'd298},{  1'b0, 1'b0, 8'd152,  9'd277},{  1'b0, 1'b0, 8'd148,    9'd0},{  1'b0, 1'b0, 8'd134,  9'd194},{  1'b0, 1'b0, 8'd130,    9'd0},{  1'b0, 1'b0, 8'd126,  9'd324},{  1'b0, 1'b0, 8'd115,  9'd223},{  1'b0, 1'b0, 8'd114,  9'd180},{  1'b0, 1'b0, 8'd112,    9'd0},{  1'b0, 1'b0,  8'd94,    9'd0},{  1'b0, 1'b0,  8'd90,   9'd98},{  1'b0, 1'b0,  8'd90,  9'd180},{  1'b0, 1'b0,  8'd80,  9'd129},{  1'b0, 1'b0,  8'd77,  9'd161},{  1'b0, 1'b0,  8'd76,    9'd0},{  1'b0, 1'b0,  8'd68,  9'd246},{  1'b0, 1'b0,  8'd61,   9'd65},{  1'b0, 1'b0,  8'd58,    9'd0},{  1'b0, 1'b0,  8'd51,  9'd128},{  1'b0, 1'b0,  8'd45,   9'd33},{  1'b0, 1'b0,  8'd40,    9'd0},{  1'b0, 1'b0,  8'd24,  9'd159},{  1'b0, 1'b0,  8'd22,    9'd0},{  1'b0, 1'b0,  8'd22,   9'd75},{  1'b0, 1'b0,  8'd14,   9'd82},{  1'b0, 1'b0,   8'd5,  9'd121},{  1'b0, 1'b0,   8'd4,    9'd0},{  1'b0, 1'b1,   8'd4,  9'd313},
{  1'b0, 1'b0, 8'd167,    9'd0},{  1'b0, 1'b0, 8'd166,    9'd0},{  1'b0, 1'b0, 8'd159,  9'd149},{  1'b0, 1'b0, 8'd149,    9'd0},{  1'b0, 1'b0, 8'd149,   9'd84},{  1'b0, 1'b0, 8'd133,  9'd311},{  1'b0, 1'b0, 8'd132,  9'd351},{  1'b0, 1'b0, 8'd131,    9'd0},{  1'b0, 1'b0, 8'd122,  9'd173},{  1'b0, 1'b0, 8'd121,  9'd211},{  1'b0, 1'b0, 8'd113,    9'd0},{  1'b0, 1'b0, 8'd105,   9'd16},{  1'b0, 1'b0,  8'd95,    9'd0},{  1'b0, 1'b0,  8'd92,   9'd88},{  1'b0, 1'b0,  8'd77,    9'd0},{  1'b0, 1'b0,  8'd74,  9'd246},{  1'b0, 1'b0,  8'd74,  9'd242},{  1'b0, 1'b0,  8'd61,    9'd7},{  1'b0, 1'b0,  8'd59,    9'd0},{  1'b0, 1'b0,  8'd59,  9'd307},{  1'b0, 1'b0,  8'd46,  9'd300},{  1'b0, 1'b0,  8'd46,   9'd26},{  1'b0, 1'b0,  8'd41,    9'd0},{  1'b0, 1'b0,  8'd32,  9'd238},{  1'b0, 1'b0,  8'd23,    9'd0},{  1'b0, 1'b0,  8'd18,  9'd300},{  1'b0, 1'b0,  8'd16,  9'd231},{  1'b0, 1'b0,  8'd11,  9'd164},{  1'b0, 1'b0,   8'd8,  9'd145},{  1'b0, 1'b1,   8'd5,    9'd0},
{  1'b0, 1'b0, 8'd168,    9'd0},{  1'b0, 1'b0, 8'd167,    9'd0},{  1'b0, 1'b0, 8'd151,  9'd293},{  1'b0, 1'b0, 8'd150,    9'd0},{  1'b0, 1'b0, 8'd148,  9'd214},{  1'b0, 1'b0, 8'd139,  9'd145},{  1'b0, 1'b0, 8'd135,  9'd195},{  1'b0, 1'b0, 8'd132,    9'd0},{  1'b0, 1'b0, 8'd121,  9'd279},{  1'b0, 1'b0, 8'd114,    9'd0},{  1'b0, 1'b0, 8'd113,  9'd145},{  1'b0, 1'b0,  8'd96,    9'd0},{  1'b0, 1'b0,  8'd95,  9'd150},{  1'b0, 1'b0,  8'd93,  9'd286},{  1'b0, 1'b0,  8'd87,  9'd319},{  1'b0, 1'b0,  8'd78,    9'd0},{  1'b0, 1'b0,  8'd78,  9'd151},{  1'b0, 1'b0,  8'd68,   9'd50},{  1'b0, 1'b0,  8'd60,    9'd0},{  1'b0, 1'b0,  8'd60,  9'd253},{  1'b0, 1'b0,  8'd52,   9'd62},{  1'b0, 1'b0,  8'd42,    9'd0},{  1'b0, 1'b0,  8'd40,  9'd197},{  1'b0, 1'b0,  8'd24,    9'd0},{  1'b0, 1'b0,  8'd21,  9'd308},{  1'b0, 1'b0,  8'd19,  9'd166},{  1'b0, 1'b0,   8'd8,  9'd296},{  1'b0, 1'b0,   8'd6,    9'd0},{  1'b0, 1'b0,   8'd5,   9'd96},{  1'b0, 1'b1,   8'd2,   9'd46},
{  1'b0, 1'b0, 8'd169,    9'd0},{  1'b0, 1'b0, 8'd168,    9'd0},{  1'b0, 1'b0, 8'd156,   9'd78},{  1'b0, 1'b0, 8'd151,    9'd0},{  1'b0, 1'b0, 8'd148,  9'd286},{  1'b0, 1'b0, 8'd136,  9'd127},{  1'b0, 1'b0, 8'd134,   9'd72},{  1'b0, 1'b0, 8'd133,    9'd0},{  1'b0, 1'b0, 8'd116,  9'd125},{  1'b0, 1'b0, 8'd116,  9'd170},{  1'b0, 1'b0, 8'd115,    9'd0},{  1'b0, 1'b0,  8'd97,    9'd0},{  1'b0, 1'b0,  8'd92,  9'd238},{  1'b0, 1'b0,  8'd91,  9'd119},{  1'b0, 1'b0,  8'd84,  9'd342},{  1'b0, 1'b0,  8'd81,  9'd311},{  1'b0, 1'b0,  8'd79,    9'd0},{  1'b0, 1'b0,  8'd61,    9'd0},{  1'b0, 1'b0,  8'd58,  9'd195},{  1'b0, 1'b0,  8'd56,   9'd68},{  1'b0, 1'b0,  8'd43,    9'd0},{  1'b0, 1'b0,  8'd41,  9'd306},{  1'b0, 1'b0,  8'd36,  9'd231},{  1'b0, 1'b0,  8'd28,  9'd273},{  1'b0, 1'b0,  8'd25,    9'd0},{  1'b0, 1'b0,  8'd24,  9'd301},{  1'b0, 1'b0,   8'd7,    9'd0},{  1'b0, 1'b0,   8'd7,  9'd121},{  1'b0, 1'b0,   8'd1,  9'd267},{  1'b0, 1'b1,   8'd0,  9'd142},
{  1'b0, 1'b0, 8'd170,    9'd0},{  1'b0, 1'b0, 8'd169,    9'd0},{  1'b0, 1'b0, 8'd161,  9'd188},{  1'b0, 1'b0, 8'd152,    9'd0},{  1'b0, 1'b0, 8'd150,  9'd175},{  1'b0, 1'b0, 8'd141,  9'd346},{  1'b0, 1'b0, 8'd134,    9'd0},{  1'b0, 1'b0, 8'd131,   9'd82},{  1'b0, 1'b0, 8'd118,   9'd66},{  1'b0, 1'b0, 8'd116,    9'd0},{  1'b0, 1'b0, 8'd109,  9'd117},{  1'b0, 1'b0, 8'd107,  9'd354},{  1'b0, 1'b0, 8'd102,  9'd341},{  1'b0, 1'b0,  8'd98,    9'd0},{  1'b0, 1'b0,  8'd88,  9'd336},{  1'b0, 1'b0,  8'd88,  9'd181},{  1'b0, 1'b0,  8'd80,    9'd0},{  1'b0, 1'b0,  8'd63,   9'd60},{  1'b0, 1'b0,  8'd62,    9'd0},{  1'b0, 1'b0,  8'd55,   9'd43},{  1'b0, 1'b0,  8'd47,  9'd262},{  1'b0, 1'b0,  8'd47,  9'd289},{  1'b0, 1'b0,  8'd44,    9'd0},{  1'b0, 1'b0,  8'd30,   9'd79},{  1'b0, 1'b0,  8'd26,    9'd0},{  1'b0, 1'b0,  8'd26,  9'd143},{  1'b0, 1'b0,  8'd17,   9'd14},{  1'b0, 1'b0,  8'd11,  9'd243},{  1'b0, 1'b0,   8'd8,    9'd0},{  1'b0, 1'b1,   8'd6,  9'd315},
{  1'b0, 1'b0, 8'd171,    9'd0},{  1'b0, 1'b0, 8'd170,    9'd0},{  1'b0, 1'b0, 8'd160,   9'd97},{  1'b0, 1'b0, 8'd153,    9'd0},{  1'b0, 1'b0, 8'd145,  9'd133},{  1'b0, 1'b0, 8'd140,  9'd181},{  1'b0, 1'b0, 8'd135,    9'd0},{  1'b0, 1'b0, 8'd128,  9'd342},{  1'b0, 1'b0, 8'd123,  9'd265},{  1'b0, 1'b0, 8'd120,  9'd254},{  1'b0, 1'b0, 8'd117,    9'd0},{  1'b0, 1'b0, 8'd106,  9'd330},{  1'b0, 1'b0,  8'd99,    9'd0},{  1'b0, 1'b0,  8'd97,   9'd38},{  1'b0, 1'b0,  8'd81,    9'd0},{  1'b0, 1'b0,  8'd80,  9'd333},{  1'b0, 1'b0,  8'd72,   9'd47},{  1'b0, 1'b0,  8'd70,  9'd143},{  1'b0, 1'b0,  8'd63,    9'd0},{  1'b0, 1'b0,  8'd60,  9'd107},{  1'b0, 1'b0,  8'd45,    9'd0},{  1'b0, 1'b0,  8'd43,   9'd42},{  1'b0, 1'b0,  8'd42,   9'd95},{  1'b0, 1'b0,  8'd27,    9'd0},{  1'b0, 1'b0,  8'd27,   9'd65},{  1'b0, 1'b0,  8'd23,    9'd6},{  1'b0, 1'b0,  8'd15,  9'd213},{  1'b0, 1'b0,   8'd9,    9'd0},{  1'b0, 1'b0,   8'd9,   9'd97},{  1'b0, 1'b1,   8'd2,    9'd4},
{  1'b0, 1'b0, 8'd172,    9'd0},{  1'b0, 1'b0, 8'd171,    9'd0},{  1'b0, 1'b0, 8'd160,   9'd17},{  1'b0, 1'b0, 8'd154,    9'd0},{  1'b0, 1'b0, 8'd154,  9'd242},{  1'b0, 1'b0, 8'd139,  9'd156},{  1'b0, 1'b0, 8'd136,    9'd0},{  1'b0, 1'b0, 8'd132,  9'd224},{  1'b0, 1'b0, 8'd118,    9'd0},{  1'b0, 1'b0, 8'd114,   9'd56},{  1'b0, 1'b0, 8'd108,  9'd260},{  1'b0, 1'b0, 8'd104,  9'd285},{  1'b0, 1'b0, 8'd100,    9'd0},{  1'b0, 1'b0,  8'd93,   9'd69},{  1'b0, 1'b0,  8'd89,  9'd184},{  1'b0, 1'b0,  8'd82,    9'd0},{  1'b0, 1'b0,  8'd73,  9'd220},{  1'b0, 1'b0,  8'd67,  9'd154},{  1'b0, 1'b0,  8'd64,    9'd0},{  1'b0, 1'b0,  8'd54,  9'd326},{  1'b0, 1'b0,  8'd51,  9'd171},{  1'b0, 1'b0,  8'd46,    9'd0},{  1'b0, 1'b0,  8'd38,   9'd48},{  1'b0, 1'b0,  8'd33,  9'd298},{  1'b0, 1'b0,  8'd32,  9'd102},{  1'b0, 1'b0,  8'd28,    9'd0},{  1'b0, 1'b0,  8'd17,  9'd131},{  1'b0, 1'b0,  8'd14,   9'd59},{  1'b0, 1'b0,  8'd10,    9'd0},{  1'b0, 1'b1,  8'd10,  9'd174},
{  1'b0, 1'b0, 8'd173,    9'd0},{  1'b0, 1'b0, 8'd172,    9'd0},{  1'b0, 1'b0, 8'd161,  9'd110},{  1'b0, 1'b0, 8'd155,    9'd0},{  1'b0, 1'b0, 8'd147,  9'd311},{  1'b0, 1'b0, 8'd137,    9'd0},{  1'b0, 1'b0, 8'd137,  9'd213},{  1'b0, 1'b0, 8'd130,  9'd123},{  1'b0, 1'b0, 8'd120,  9'd210},{  1'b0, 1'b0, 8'd119,    9'd0},{  1'b0, 1'b0, 8'd111,   9'd97},{  1'b0, 1'b0, 8'd102,  9'd184},{  1'b0, 1'b0, 8'd101,    9'd0},{  1'b0, 1'b0, 8'd101,  9'd284},{  1'b0, 1'b0,  8'd83,    9'd0},{  1'b0, 1'b0,  8'd73,  9'd227},{  1'b0, 1'b0,  8'd72,  9'd248},{  1'b0, 1'b0,  8'd67,   9'd10},{  1'b0, 1'b0,  8'd65,    9'd0},{  1'b0, 1'b0,  8'd55,  9'd186},{  1'b0, 1'b0,  8'd48,    9'd8},{  1'b0, 1'b0,  8'd47,    9'd0},{  1'b0, 1'b0,  8'd38,  9'd155},{  1'b0, 1'b0,  8'd34,   9'd98},{  1'b0, 1'b0,  8'd29,    9'd0},{  1'b0, 1'b0,  8'd29,  9'd125},{  1'b0, 1'b0,  8'd12,  9'd176},{  1'b0, 1'b0,  8'd11,    9'd0},{  1'b0, 1'b0,   8'd4,   9'd58},{  1'b0, 1'b1,   8'd1,  9'd174},
{  1'b0, 1'b0, 8'd174,    9'd0},{  1'b0, 1'b0, 8'd173,    9'd0},{  1'b0, 1'b0, 8'd158,   9'd85},{  1'b0, 1'b0, 8'd156,    9'd0},{  1'b0, 1'b0, 8'd144,   9'd88},{  1'b0, 1'b0, 8'd138,    9'd0},{  1'b0, 1'b0, 8'd130,  9'd352},{  1'b0, 1'b0, 8'd129,  9'd196},{  1'b0, 1'b0, 8'd120,    9'd0},{  1'b0, 1'b0, 8'd119,  9'd217},{  1'b0, 1'b0, 8'd110,  9'd354},{  1'b0, 1'b0, 8'd107,  9'd252},{  1'b0, 1'b0, 8'd102,    9'd0},{  1'b0, 1'b0,  8'd96,  9'd186},{  1'b0, 1'b0,  8'd84,    9'd0},{  1'b0, 1'b0,  8'd83,   9'd54},{  1'b0, 1'b0,  8'd76,   9'd63},{  1'b0, 1'b0,  8'd66,    9'd0},{  1'b0, 1'b0,  8'd66,  9'd196},{  1'b0, 1'b0,  8'd64,  9'd246},{  1'b0, 1'b0,  8'd50,   9'd64},{  1'b0, 1'b0,  8'd48,    9'd0},{  1'b0, 1'b0,  8'd42,   9'd28},{  1'b0, 1'b0,  8'd35,  9'd178},{  1'b0, 1'b0,  8'd31,   9'd26},{  1'b0, 1'b0,  8'd30,    9'd0},{  1'b0, 1'b0,  8'd12,    9'd0},{  1'b0, 1'b0,   8'd9,  9'd213},{  1'b0, 1'b0,   8'd7,   9'd30},{  1'b0, 1'b1,   8'd6,  9'd185},
{  1'b0, 1'b0, 8'd175,    9'd0},{  1'b0, 1'b0, 8'd174,    9'd0},{  1'b0, 1'b0, 8'd157,    9'd0},{  1'b0, 1'b0, 8'd157,  9'd313},{  1'b0, 1'b0, 8'd145,   9'd68},{  1'b0, 1'b0, 8'd139,    9'd0},{  1'b0, 1'b0, 8'd138,   9'd35},{  1'b0, 1'b0, 8'd136,  9'd286},{  1'b0, 1'b0, 8'd125,  9'd243},{  1'b0, 1'b0, 8'd121,    9'd0},{  1'b0, 1'b0, 8'd117,  9'd170},{  1'b0, 1'b0, 8'd103,    9'd0},{  1'b0, 1'b0, 8'd103,  9'd107},{  1'b0, 1'b0, 8'd101,   9'd51},{  1'b0, 1'b0,  8'd85,    9'd0},{  1'b0, 1'b0,  8'd85,  9'd297},{  1'b0, 1'b0,  8'd82,   9'd87},{  1'b0, 1'b0,  8'd69,   9'd61},{  1'b0, 1'b0,  8'd67,    9'd0},{  1'b0, 1'b0,  8'd57,  9'd234},{  1'b0, 1'b0,  8'd49,    9'd0},{  1'b0, 1'b0,  8'd45,  9'd312},{  1'b0, 1'b0,  8'd43,  9'd201},{  1'b0, 1'b0,  8'd31,    9'd0},{  1'b0, 1'b0,  8'd29,  9'd330},{  1'b0, 1'b0,  8'd20,   9'd92},{  1'b0, 1'b0,  8'd15,   9'd98},{  1'b0, 1'b0,  8'd15,  9'd242},{  1'b0, 1'b0,  8'd13,    9'd0},{  1'b0, 1'b1,   8'd0,  9'd311},
{  1'b0, 1'b0, 8'd176,    9'd0},{  1'b0, 1'b0, 8'd175,    9'd0},{  1'b0, 1'b0, 8'd158,    9'd0},{  1'b0, 1'b0, 8'd153,  9'd313},{  1'b0, 1'b0, 8'd147,   9'd39},{  1'b0, 1'b0, 8'd142,  9'd163},{  1'b0, 1'b0, 8'd140,    9'd0},{  1'b0, 1'b0, 8'd127,  9'd284},{  1'b0, 1'b0, 8'd122,    9'd0},{  1'b0, 1'b0, 8'd122,  9'd194},{  1'b0, 1'b0, 8'd113,   9'd66},{  1'b0, 1'b0, 8'd104,    9'd0},{  1'b0, 1'b0,  8'd99,   9'd41},{  1'b0, 1'b0,  8'd95,  9'd267},{  1'b0, 1'b0,  8'd86,    9'd0},{  1'b0, 1'b0,  8'd81,  9'd332},{  1'b0, 1'b0,  8'd75,  9'd288},{  1'b0, 1'b0,  8'd70,  9'd349},{  1'b0, 1'b0,  8'd68,    9'd0},{  1'b0, 1'b0,  8'd65,  9'd237},{  1'b0, 1'b0,  8'd50,    9'd0},{  1'b0, 1'b0,  8'd48,  9'd101},{  1'b0, 1'b0,  8'd41,  9'd159},{  1'b0, 1'b0,  8'd32,    9'd0},{  1'b0, 1'b0,  8'd21,  9'd257},{  1'b0, 1'b0,  8'd19,  9'd242},{  1'b0, 1'b0,  8'd14,    9'd0},{  1'b0, 1'b0,  8'd10,  9'd230},{  1'b0, 1'b0,   8'd6,  9'd124},{  1'b0, 1'b1,   8'd3,  9'd225},
{  1'b0, 1'b0, 8'd177,    9'd0},{  1'b0, 1'b0, 8'd176,    9'd0},{  1'b0, 1'b0, 8'd159,    9'd0},{  1'b0, 1'b0, 8'd155,  9'd197},{  1'b0, 1'b0, 8'd151,  9'd146},{  1'b0, 1'b0, 8'd141,    9'd0},{  1'b0, 1'b0, 8'd129,  9'd138},{  1'b0, 1'b0, 8'd128,  9'd317},{  1'b0, 1'b0, 8'd123,    9'd0},{  1'b0, 1'b0, 8'd115,  9'd293},{  1'b0, 1'b0, 8'd112,  9'd155},{  1'b0, 1'b0, 8'd105,    9'd0},{  1'b0, 1'b0, 8'd104,   9'd79},{  1'b0, 1'b0,  8'd99,  9'd116},{  1'b0, 1'b0,  8'd87,    9'd0},{  1'b0, 1'b0,  8'd85,  9'd220},{  1'b0, 1'b0,  8'd83,  9'd244},{  1'b0, 1'b0,  8'd69,    9'd0},{  1'b0, 1'b0,  8'd66,   9'd20},{  1'b0, 1'b0,  8'd63,  9'd173},{  1'b0, 1'b0,  8'd51,    9'd0},{  1'b0, 1'b0,  8'd49,   9'd93},{  1'b0, 1'b0,  8'd49,  9'd123},{  1'b0, 1'b0,  8'd33,    9'd0},{  1'b0, 1'b0,  8'd28,   9'd51},{  1'b0, 1'b0,  8'd22,  9'd217},{  1'b0, 1'b0,  8'd17,  9'd280},{  1'b0, 1'b0,  8'd15,    9'd0},{  1'b0, 1'b0,  8'd13,  9'd336},{  1'b0, 1'b1,   8'd2,  9'd137},
{  1'b0, 1'b0, 8'd178,    9'd0},{  1'b0, 1'b0, 8'd177,    9'd0},{  1'b0, 1'b0, 8'd160,    9'd0},{  1'b0, 1'b0, 8'd150,  9'd141},{  1'b0, 1'b0, 8'd149,   9'd72},{  1'b0, 1'b0, 8'd142,    9'd0},{  1'b0, 1'b0, 8'd142,   9'd35},{  1'b0, 1'b0, 8'd127,   9'd59},{  1'b0, 1'b0, 8'd125,  9'd226},{  1'b0, 1'b0, 8'd124,    9'd0},{  1'b0, 1'b0, 8'd111,  9'd317},{  1'b0, 1'b0, 8'd106,    9'd0},{  1'b0, 1'b0, 8'd103,  9'd277},{  1'b0, 1'b0,  8'd98,  9'd230},{  1'b0, 1'b0,  8'd88,    9'd0},{  1'b0, 1'b0,  8'd77,  9'd177},{  1'b0, 1'b0,  8'd76,  9'd245},{  1'b0, 1'b0,  8'd70,    9'd0},{  1'b0, 1'b0,  8'd65,  9'd317},{  1'b0, 1'b0,  8'd59,  9'd176},{  1'b0, 1'b0,  8'd53,  9'd319},{  1'b0, 1'b0,  8'd52,    9'd0},{  1'b0, 1'b0,  8'd37,  9'd160},{  1'b0, 1'b0,  8'd34,    9'd0},{  1'b0, 1'b0,  8'd33,  9'd344},{  1'b0, 1'b0,  8'd18,  9'd339},{  1'b0, 1'b0,  8'd16,    9'd0},{  1'b0, 1'b0,  8'd14,  9'd299},{  1'b0, 1'b0,   8'd9,   9'd85},{  1'b0, 1'b1,   8'd4,  9'd161},
{  1'b0, 1'b0, 8'd179,    9'd0},{  1'b0, 1'b0, 8'd178,    9'd0},{  1'b0, 1'b0, 8'd161,    9'd0},{  1'b0, 1'b0, 8'd157,  9'd258},{  1'b0, 1'b0, 8'd156,  9'd198},{  1'b0, 1'b0, 8'd143,    9'd0},{  1'b0, 1'b0, 8'd141,   9'd32},{  1'b0, 1'b0, 8'd133,   9'd72},{  1'b0, 1'b0, 8'd125,    9'd0},{  1'b0, 1'b0, 8'd123,   9'd23},{  1'b0, 1'b0, 8'd117,  9'd137},{  1'b0, 1'b0, 8'd107,    9'd0},{  1'b0, 1'b0,  8'd96,   9'd81},{  1'b0, 1'b0,  8'd94,  9'd329},{  1'b0, 1'b0,  8'd89,    9'd0},{  1'b0, 1'b0,  8'd89,  9'd226},{  1'b0, 1'b0,  8'd86,  9'd105},{  1'b0, 1'b0,  8'd71,    9'd0},{  1'b0, 1'b0,  8'd71,   9'd80},{  1'b0, 1'b0,  8'd54,  9'd144},{  1'b0, 1'b0,  8'd53,    9'd0},{  1'b0, 1'b0,  8'd50,   9'd24},{  1'b0, 1'b0,  8'd39,  9'd309},{  1'b0, 1'b0,  8'd35,    9'd0},{  1'b0, 1'b0,  8'd25,  9'd335},{  1'b0, 1'b0,  8'd25,   9'd37},{  1'b0, 1'b0,  8'd17,    9'd0},{  1'b0, 1'b0,  8'd13,   9'd78},{  1'b0, 1'b0,  8'd10,  9'd308},{  1'b0, 1'b1,   8'd3,  9'd236}
};
localparam bit [18 : 0] cLARGE_HS_V_TAB_9BY10_PACKED[cLARGE_HS_TAB_9BY10_PACKED_SIZE] = '{
{8'd179, 1'b0,   10'd0},{8'd179, 1'b1, 10'd510},
{8'd178, 1'b0, 10'd480},{8'd178, 1'b1, 10'd511},
{8'd177, 1'b0, 10'd450},{8'd177, 1'b1, 10'd481},
{8'd176, 1'b0, 10'd420},{8'd176, 1'b1, 10'd451},
{8'd175, 1'b0, 10'd390},{8'd175, 1'b1, 10'd421},
{8'd174, 1'b0, 10'd360},{8'd174, 1'b1, 10'd391},
{8'd173, 1'b0, 10'd330},{8'd173, 1'b1, 10'd361},
{8'd172, 1'b0, 10'd300},{8'd172, 1'b1, 10'd331},
{8'd171, 1'b0, 10'd270},{8'd171, 1'b1, 10'd301},
{8'd170, 1'b0, 10'd240},{8'd170, 1'b1, 10'd271},
{8'd169, 1'b0, 10'd210},{8'd169, 1'b1, 10'd241},
{8'd168, 1'b0, 10'd180},{8'd168, 1'b1, 10'd211},
{8'd167, 1'b0, 10'd150},{8'd167, 1'b1, 10'd181},
{8'd166, 1'b0, 10'd120},{8'd166, 1'b1, 10'd151},
{8'd165, 1'b0,  10'd90},{8'd165, 1'b1, 10'd121},
{8'd164, 1'b0,  10'd60},{8'd164, 1'b1,  10'd91},
{8'd163, 1'b0,  10'd30},{8'd163, 1'b1,  10'd61},
{8'd162, 1'b0,   10'd1},{8'd162, 1'b1,  10'd31},
{8'd161, 1'b0, 10'd242},{8'd161, 1'b0, 10'd332},{8'd161, 1'b1, 10'd512},
{8'd160, 1'b0, 10'd272},{8'd160, 1'b0, 10'd302},{8'd160, 1'b1, 10'd482},
{8'd159, 1'b0,  10'd62},{8'd159, 1'b0, 10'd152},{8'd159, 1'b1, 10'd452},
{8'd158, 1'b0,  10'd32},{8'd158, 1'b0, 10'd362},{8'd158, 1'b1, 10'd422},
{8'd157, 1'b0, 10'd392},{8'd157, 1'b0, 10'd393},{8'd157, 1'b1, 10'd513},
{8'd156, 1'b0, 10'd212},{8'd156, 1'b0, 10'd363},{8'd156, 1'b1, 10'd514},
{8'd155, 1'b0, 10'd122},{8'd155, 1'b0, 10'd333},{8'd155, 1'b1, 10'd453},
{8'd154, 1'b0,   10'd2},{8'd154, 1'b0, 10'd303},{8'd154, 1'b1, 10'd304},
{8'd153, 1'b0,   10'd3},{8'd153, 1'b0, 10'd273},{8'd153, 1'b1, 10'd423},
{8'd152, 1'b0,  10'd92},{8'd152, 1'b0, 10'd123},{8'd152, 1'b1, 10'd243},
{8'd151, 1'b0, 10'd182},{8'd151, 1'b0, 10'd213},{8'd151, 1'b1, 10'd454},
{8'd150, 1'b0, 10'd183},{8'd150, 1'b0, 10'd244},{8'd150, 1'b1, 10'd483},
{8'd149, 1'b0, 10'd153},{8'd149, 1'b0, 10'd154},{8'd149, 1'b1, 10'd484},
{8'd148, 1'b0, 10'd124},{8'd148, 1'b0, 10'd184},{8'd148, 1'b1, 10'd214},
{8'd147, 1'b0,  10'd93},{8'd147, 1'b0, 10'd334},{8'd147, 1'b1, 10'd424},
{8'd146, 1'b0,  10'd63},{8'd146, 1'b0,  10'd64},{8'd146, 1'b1,  10'd94},
{8'd145, 1'b0,  10'd33},{8'd145, 1'b0, 10'd274},{8'd145, 1'b1, 10'd394},
{8'd144, 1'b0,   10'd4},{8'd144, 1'b0,  10'd34},{8'd144, 1'b1, 10'd364},
{8'd143, 1'b0,  10'd35},{8'd143, 1'b0,  10'd65},{8'd143, 1'b1, 10'd515},
{8'd142, 1'b0, 10'd425},{8'd142, 1'b0, 10'd485},{8'd142, 1'b1, 10'd486},
{8'd141, 1'b0, 10'd245},{8'd141, 1'b0, 10'd455},{8'd141, 1'b1, 10'd516},
{8'd140, 1'b0,  10'd36},{8'd140, 1'b0, 10'd275},{8'd140, 1'b1, 10'd426},
{8'd139, 1'b0, 10'd185},{8'd139, 1'b0, 10'd305},{8'd139, 1'b1, 10'd395},
{8'd138, 1'b0,  10'd95},{8'd138, 1'b0, 10'd365},{8'd138, 1'b1, 10'd396},
{8'd137, 1'b0,  10'd66},{8'd137, 1'b0, 10'd335},{8'd137, 1'b1, 10'd336},
{8'd136, 1'b0, 10'd215},{8'd136, 1'b0, 10'd306},{8'd136, 1'b1, 10'd397},
{8'd135, 1'b0,  10'd96},{8'd135, 1'b0, 10'd186},{8'd135, 1'b1, 10'd276},
{8'd134, 1'b0, 10'd125},{8'd134, 1'b0, 10'd216},{8'd134, 1'b1, 10'd246},
{8'd133, 1'b0, 10'd155},{8'd133, 1'b0, 10'd217},{8'd133, 1'b1, 10'd517},
{8'd132, 1'b0, 10'd156},{8'd132, 1'b0, 10'd187},{8'd132, 1'b1, 10'd307},
{8'd131, 1'b0,   10'd5},{8'd131, 1'b0, 10'd157},{8'd131, 1'b1, 10'd247},
{8'd130, 1'b0, 10'd126},{8'd130, 1'b0, 10'd337},{8'd130, 1'b1, 10'd366},
{8'd129, 1'b0,  10'd97},{8'd129, 1'b0, 10'd367},{8'd129, 1'b1, 10'd456},
{8'd128, 1'b0,  10'd67},{8'd128, 1'b0, 10'd277},{8'd128, 1'b1, 10'd457},
{8'd127, 1'b0,  10'd37},{8'd127, 1'b0, 10'd427},{8'd127, 1'b1, 10'd487},
{8'd126, 1'b0,   10'd6},{8'd126, 1'b0,   10'd7},{8'd126, 1'b1, 10'd127},
{8'd125, 1'b0, 10'd398},{8'd125, 1'b0, 10'd488},{8'd125, 1'b1, 10'd518},
{8'd124, 1'b0,   10'd8},{8'd124, 1'b0,  10'd68},{8'd124, 1'b1, 10'd489},
{8'd123, 1'b0, 10'd278},{8'd123, 1'b0, 10'd458},{8'd123, 1'b1, 10'd519},
{8'd122, 1'b0, 10'd158},{8'd122, 1'b0, 10'd428},{8'd122, 1'b1, 10'd429},
{8'd121, 1'b0, 10'd159},{8'd121, 1'b0, 10'd188},{8'd121, 1'b1, 10'd399},
{8'd120, 1'b0, 10'd279},{8'd120, 1'b0, 10'd338},{8'd120, 1'b1, 10'd368},
{8'd119, 1'b0,  10'd38},{8'd119, 1'b0, 10'd339},{8'd119, 1'b1, 10'd369},
{8'd118, 1'b0,  10'd39},{8'd118, 1'b0, 10'd248},{8'd118, 1'b1, 10'd308},
{8'd117, 1'b0, 10'd280},{8'd117, 1'b0, 10'd400},{8'd117, 1'b1, 10'd520},
{8'd116, 1'b0, 10'd218},{8'd116, 1'b0, 10'd219},{8'd116, 1'b1, 10'd249},
{8'd115, 1'b0, 10'd128},{8'd115, 1'b0, 10'd220},{8'd115, 1'b1, 10'd459},
{8'd114, 1'b0, 10'd129},{8'd114, 1'b0, 10'd189},{8'd114, 1'b1, 10'd309},
{8'd113, 1'b0, 10'd160},{8'd113, 1'b0, 10'd190},{8'd113, 1'b1, 10'd430},
{8'd112, 1'b0,   10'd9},{8'd112, 1'b0, 10'd130},{8'd112, 1'b1, 10'd460},
{8'd111, 1'b0,  10'd98},{8'd111, 1'b0, 10'd340},{8'd111, 1'b1, 10'd490},
{8'd110, 1'b0,  10'd69},{8'd110, 1'b0,  10'd99},{8'd110, 1'b1, 10'd370},
{8'd109, 1'b0,  10'd40},{8'd109, 1'b0,  10'd70},{8'd109, 1'b1, 10'd250},
{8'd108, 1'b0,  10'd10},{8'd108, 1'b0, 10'd100},{8'd108, 1'b1, 10'd310},
{8'd107, 1'b0, 10'd251},{8'd107, 1'b0, 10'd371},{8'd107, 1'b1, 10'd521},
{8'd106, 1'b0, 10'd101},{8'd106, 1'b0, 10'd281},{8'd106, 1'b1, 10'd491},
{8'd105, 1'b0, 10'd102},{8'd105, 1'b0, 10'd161},{8'd105, 1'b1, 10'd461},
{8'd104, 1'b0, 10'd311},{8'd104, 1'b0, 10'd431},{8'd104, 1'b1, 10'd462},
{8'd103, 1'b0, 10'd401},{8'd103, 1'b0, 10'd402},{8'd103, 1'b1, 10'd492},
{8'd102, 1'b0, 10'd252},{8'd102, 1'b0, 10'd341},{8'd102, 1'b1, 10'd372},
{8'd101, 1'b0, 10'd342},{8'd101, 1'b0, 10'd343},{8'd101, 1'b1, 10'd403},
{8'd100, 1'b0,  10'd41},{8'd100, 1'b0,  10'd71},{8'd100, 1'b1, 10'd312},
{ 8'd99, 1'b0, 10'd282},{ 8'd99, 1'b0, 10'd432},{ 8'd99, 1'b1, 10'd463},
{ 8'd98, 1'b0,  10'd72},{ 8'd98, 1'b0, 10'd253},{ 8'd98, 1'b1, 10'd493},
{ 8'd97, 1'b0,  10'd11},{ 8'd97, 1'b0, 10'd221},{ 8'd97, 1'b1, 10'd283},
{ 8'd96, 1'b0, 10'd191},{ 8'd96, 1'b0, 10'd373},{ 8'd96, 1'b1, 10'd522},
{ 8'd95, 1'b0, 10'd162},{ 8'd95, 1'b0, 10'd192},{ 8'd95, 1'b1, 10'd433},
{ 8'd94, 1'b0,  10'd42},{ 8'd94, 1'b0, 10'd131},{ 8'd94, 1'b1, 10'd523},
{ 8'd93, 1'b0, 10'd103},{ 8'd93, 1'b0, 10'd193},{ 8'd93, 1'b1, 10'd313},
{ 8'd92, 1'b0,  10'd73},{ 8'd92, 1'b0, 10'd163},{ 8'd92, 1'b1, 10'd222},
{ 8'd91, 1'b0,  10'd12},{ 8'd91, 1'b0,  10'd43},{ 8'd91, 1'b1, 10'd223},
{ 8'd90, 1'b0,  10'd13},{ 8'd90, 1'b0, 10'd132},{ 8'd90, 1'b1, 10'd133},
{ 8'd89, 1'b0, 10'd314},{ 8'd89, 1'b0, 10'd524},{ 8'd89, 1'b1, 10'd525},
{ 8'd88, 1'b0, 10'd254},{ 8'd88, 1'b0, 10'd255},{ 8'd88, 1'b1, 10'd494},
{ 8'd87, 1'b0,  10'd44},{ 8'd87, 1'b0, 10'd194},{ 8'd87, 1'b1, 10'd464},
{ 8'd86, 1'b0,  10'd14},{ 8'd86, 1'b0, 10'd434},{ 8'd86, 1'b1, 10'd526},
{ 8'd85, 1'b0, 10'd404},{ 8'd85, 1'b0, 10'd405},{ 8'd85, 1'b1, 10'd465},
{ 8'd84, 1'b0,  10'd15},{ 8'd84, 1'b0, 10'd224},{ 8'd84, 1'b1, 10'd374},
{ 8'd83, 1'b0, 10'd344},{ 8'd83, 1'b0, 10'd375},{ 8'd83, 1'b1, 10'd466},
{ 8'd82, 1'b0,  10'd74},{ 8'd82, 1'b0, 10'd315},{ 8'd82, 1'b1, 10'd406},
{ 8'd81, 1'b0, 10'd225},{ 8'd81, 1'b0, 10'd284},{ 8'd81, 1'b1, 10'd435},
{ 8'd80, 1'b0, 10'd134},{ 8'd80, 1'b0, 10'd256},{ 8'd80, 1'b1, 10'd285},
{ 8'd79, 1'b0,  10'd75},{ 8'd79, 1'b0, 10'd104},{ 8'd79, 1'b1, 10'd226},
{ 8'd78, 1'b0, 10'd105},{ 8'd78, 1'b0, 10'd195},{ 8'd78, 1'b1, 10'd196},
{ 8'd77, 1'b0, 10'd135},{ 8'd77, 1'b0, 10'd164},{ 8'd77, 1'b1, 10'd495},
{ 8'd76, 1'b0, 10'd136},{ 8'd76, 1'b0, 10'd376},{ 8'd76, 1'b1, 10'd496},
{ 8'd75, 1'b0,  10'd45},{ 8'd75, 1'b0, 10'd106},{ 8'd75, 1'b1, 10'd436},
{ 8'd74, 1'b0,  10'd76},{ 8'd74, 1'b0, 10'd165},{ 8'd74, 1'b1, 10'd166},
{ 8'd73, 1'b0,  10'd46},{ 8'd73, 1'b0, 10'd316},{ 8'd73, 1'b1, 10'd345},
{ 8'd72, 1'b0,  10'd16},{ 8'd72, 1'b0, 10'd286},{ 8'd72, 1'b1, 10'd346},
{ 8'd71, 1'b0, 10'd107},{ 8'd71, 1'b0, 10'd527},{ 8'd71, 1'b1, 10'd528},
{ 8'd70, 1'b0, 10'd287},{ 8'd70, 1'b0, 10'd437},{ 8'd70, 1'b1, 10'd497},
{ 8'd69, 1'b0, 10'd108},{ 8'd69, 1'b0, 10'd407},{ 8'd69, 1'b1, 10'd467},
{ 8'd68, 1'b0, 10'd137},{ 8'd68, 1'b0, 10'd197},{ 8'd68, 1'b1, 10'd438},
{ 8'd67, 1'b0, 10'd317},{ 8'd67, 1'b0, 10'd347},{ 8'd67, 1'b1, 10'd408},
{ 8'd66, 1'b0, 10'd377},{ 8'd66, 1'b0, 10'd378},{ 8'd66, 1'b1, 10'd468},
{ 8'd65, 1'b0, 10'd348},{ 8'd65, 1'b0, 10'd439},{ 8'd65, 1'b1, 10'd498},
{ 8'd64, 1'b0,  10'd17},{ 8'd64, 1'b0, 10'd318},{ 8'd64, 1'b1, 10'd379},
{ 8'd63, 1'b0, 10'd257},{ 8'd63, 1'b0, 10'd288},{ 8'd63, 1'b1, 10'd469},
{ 8'd62, 1'b0,  10'd47},{ 8'd62, 1'b0,  10'd77},{ 8'd62, 1'b1, 10'd258},
{ 8'd61, 1'b0, 10'd138},{ 8'd61, 1'b0, 10'd167},{ 8'd61, 1'b1, 10'd227},
{ 8'd60, 1'b0, 10'd198},{ 8'd60, 1'b0, 10'd199},{ 8'd60, 1'b1, 10'd289},
{ 8'd59, 1'b0, 10'd168},{ 8'd59, 1'b0, 10'd169},{ 8'd59, 1'b1, 10'd499},
{ 8'd58, 1'b0,  10'd78},{ 8'd58, 1'b0, 10'd139},{ 8'd58, 1'b1, 10'd228},
{ 8'd57, 1'b0,  10'd18},{ 8'd57, 1'b0, 10'd109},{ 8'd57, 1'b1, 10'd409},
{ 8'd56, 1'b0,  10'd48},{ 8'd56, 1'b0,  10'd79},{ 8'd56, 1'b1, 10'd229},
{ 8'd55, 1'b0,  10'd49},{ 8'd55, 1'b0, 10'd259},{ 8'd55, 1'b1, 10'd349},
{ 8'd54, 1'b0,  10'd19},{ 8'd54, 1'b0, 10'd319},{ 8'd54, 1'b1, 10'd529},
{ 8'd53, 1'b0,  10'd20},{ 8'd53, 1'b0, 10'd500},{ 8'd53, 1'b1, 10'd530},
{ 8'd52, 1'b0, 10'd110},{ 8'd52, 1'b0, 10'd200},{ 8'd52, 1'b1, 10'd501},
{ 8'd51, 1'b0, 10'd140},{ 8'd51, 1'b0, 10'd320},{ 8'd51, 1'b1, 10'd470},
{ 8'd50, 1'b0, 10'd380},{ 8'd50, 1'b0, 10'd440},{ 8'd50, 1'b1, 10'd531},
{ 8'd49, 1'b0, 10'd410},{ 8'd49, 1'b0, 10'd471},{ 8'd49, 1'b1, 10'd472},
{ 8'd48, 1'b0, 10'd350},{ 8'd48, 1'b0, 10'd381},{ 8'd48, 1'b1, 10'd441},
{ 8'd47, 1'b0, 10'd260},{ 8'd47, 1'b0, 10'd261},{ 8'd47, 1'b1, 10'd351},
{ 8'd46, 1'b0, 10'd170},{ 8'd46, 1'b0, 10'd171},{ 8'd46, 1'b1, 10'd321},
{ 8'd45, 1'b0, 10'd141},{ 8'd45, 1'b0, 10'd290},{ 8'd45, 1'b1, 10'd411},
{ 8'd44, 1'b0,  10'd50},{ 8'd44, 1'b0,  10'd51},{ 8'd44, 1'b1, 10'd262},
{ 8'd43, 1'b0, 10'd230},{ 8'd43, 1'b0, 10'd291},{ 8'd43, 1'b1, 10'd412},
{ 8'd42, 1'b0, 10'd201},{ 8'd42, 1'b0, 10'd292},{ 8'd42, 1'b1, 10'd382},
{ 8'd41, 1'b0, 10'd172},{ 8'd41, 1'b0, 10'd231},{ 8'd41, 1'b1, 10'd442},
{ 8'd40, 1'b0,  10'd80},{ 8'd40, 1'b0, 10'd142},{ 8'd40, 1'b1, 10'd202},
{ 8'd39, 1'b0, 10'd111},{ 8'd39, 1'b0, 10'd112},{ 8'd39, 1'b1, 10'd532},
{ 8'd38, 1'b0,  10'd81},{ 8'd38, 1'b0, 10'd322},{ 8'd38, 1'b1, 10'd352},
{ 8'd37, 1'b0,  10'd21},{ 8'd37, 1'b0,  10'd52},{ 8'd37, 1'b1, 10'd502},
{ 8'd36, 1'b0,  10'd22},{ 8'd36, 1'b0,  10'd82},{ 8'd36, 1'b1, 10'd232},
{ 8'd35, 1'b0,  10'd23},{ 8'd35, 1'b0, 10'd383},{ 8'd35, 1'b1, 10'd533},
{ 8'd34, 1'b0,  10'd83},{ 8'd34, 1'b0, 10'd353},{ 8'd34, 1'b1, 10'd503},
{ 8'd33, 1'b0, 10'd323},{ 8'd33, 1'b0, 10'd473},{ 8'd33, 1'b1, 10'd504},
{ 8'd32, 1'b0, 10'd173},{ 8'd32, 1'b0, 10'd324},{ 8'd32, 1'b1, 10'd443},
{ 8'd31, 1'b0,  10'd53},{ 8'd31, 1'b0, 10'd384},{ 8'd31, 1'b1, 10'd413},
{ 8'd30, 1'b0,  10'd54},{ 8'd30, 1'b0, 10'd263},{ 8'd30, 1'b1, 10'd385},
{ 8'd29, 1'b0, 10'd354},{ 8'd29, 1'b0, 10'd355},{ 8'd29, 1'b1, 10'd414},
{ 8'd28, 1'b0, 10'd233},{ 8'd28, 1'b0, 10'd325},{ 8'd28, 1'b1, 10'd474},
{ 8'd27, 1'b0,  10'd84},{ 8'd27, 1'b0, 10'd293},{ 8'd27, 1'b1, 10'd294},
{ 8'd26, 1'b0,  10'd24},{ 8'd26, 1'b0, 10'd264},{ 8'd26, 1'b1, 10'd265},
{ 8'd25, 1'b0, 10'd234},{ 8'd25, 1'b0, 10'd534},{ 8'd25, 1'b1, 10'd535},
{ 8'd24, 1'b0, 10'd143},{ 8'd24, 1'b0, 10'd203},{ 8'd24, 1'b1, 10'd235},
{ 8'd23, 1'b0, 10'd113},{ 8'd23, 1'b0, 10'd174},{ 8'd23, 1'b1, 10'd295},
{ 8'd22, 1'b0, 10'd144},{ 8'd22, 1'b0, 10'd145},{ 8'd22, 1'b1, 10'd475},
{ 8'd21, 1'b0, 10'd114},{ 8'd21, 1'b0, 10'd204},{ 8'd21, 1'b1, 10'd444},
{ 8'd20, 1'b0,  10'd85},{ 8'd20, 1'b0, 10'd115},{ 8'd20, 1'b1, 10'd415},
{ 8'd19, 1'b0,  10'd55},{ 8'd19, 1'b0, 10'd205},{ 8'd19, 1'b1, 10'd445},
{ 8'd18, 1'b0,  10'd25},{ 8'd18, 1'b0, 10'd175},{ 8'd18, 1'b1, 10'd505},
{ 8'd17, 1'b0, 10'd266},{ 8'd17, 1'b0, 10'd326},{ 8'd17, 1'b0, 10'd476},{ 8'd17, 1'b1, 10'd536},
{ 8'd16, 1'b0,  10'd86},{ 8'd16, 1'b0, 10'd116},{ 8'd16, 1'b0, 10'd176},{ 8'd16, 1'b1, 10'd506},
{ 8'd15, 1'b0, 10'd296},{ 8'd15, 1'b0, 10'd416},{ 8'd15, 1'b0, 10'd417},{ 8'd15, 1'b1, 10'd477},
{ 8'd14, 1'b0, 10'd146},{ 8'd14, 1'b0, 10'd327},{ 8'd14, 1'b0, 10'd446},{ 8'd14, 1'b1, 10'd507},
{ 8'd13, 1'b0,  10'd26},{ 8'd13, 1'b0, 10'd418},{ 8'd13, 1'b0, 10'd478},{ 8'd13, 1'b1, 10'd537},
{ 8'd12, 1'b0,  10'd56},{ 8'd12, 1'b0, 10'd117},{ 8'd12, 1'b0, 10'd356},{ 8'd12, 1'b1, 10'd386},
{ 8'd11, 1'b0,  10'd27},{ 8'd11, 1'b0, 10'd177},{ 8'd11, 1'b0, 10'd267},{ 8'd11, 1'b1, 10'd357},
{ 8'd10, 1'b0, 10'd328},{ 8'd10, 1'b0, 10'd329},{ 8'd10, 1'b0, 10'd447},{ 8'd10, 1'b1, 10'd538},
{  8'd9, 1'b0, 10'd297},{  8'd9, 1'b0, 10'd298},{  8'd9, 1'b0, 10'd387},{  8'd9, 1'b1, 10'd508},
{  8'd8, 1'b0,  10'd87},{  8'd8, 1'b0, 10'd178},{  8'd8, 1'b0, 10'd206},{  8'd8, 1'b1, 10'd268},
{  8'd7, 1'b0,  10'd57},{  8'd7, 1'b0, 10'd236},{  8'd7, 1'b0, 10'd237},{  8'd7, 1'b1, 10'd388},
{  8'd6, 1'b0, 10'd207},{  8'd6, 1'b0, 10'd269},{  8'd6, 1'b0, 10'd389},{  8'd6, 1'b1, 10'd448},
{  8'd5, 1'b0, 10'd118},{  8'd5, 1'b0, 10'd147},{  8'd5, 1'b0, 10'd179},{  8'd5, 1'b1, 10'd208},
{  8'd4, 1'b0, 10'd148},{  8'd4, 1'b0, 10'd149},{  8'd4, 1'b0, 10'd358},{  8'd4, 1'b1, 10'd509},
{  8'd3, 1'b0,  10'd58},{  8'd3, 1'b0, 10'd119},{  8'd3, 1'b0, 10'd449},{  8'd3, 1'b1, 10'd539},
{  8'd2, 1'b0,  10'd88},{  8'd2, 1'b0, 10'd209},{  8'd2, 1'b0, 10'd299},{  8'd2, 1'b1, 10'd479},
{  8'd1, 1'b0,  10'd28},{  8'd1, 1'b0,  10'd59},{  8'd1, 1'b0, 10'd238},{  8'd1, 1'b1, 10'd359},
{  8'd0, 1'b0,  10'd29},{  8'd0, 1'b0,  10'd89},{  8'd0, 1'b0, 10'd239},{  8'd0, 1'b1, 10'd419}
};
