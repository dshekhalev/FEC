localparam int          cMEDIUM_HS_TAB_1BY5_PACKED_SIZE = 144;
localparam bit [17 : 0] cMEDIUM_HS_TAB_1BY5_PACKED[cMEDIUM_HS_TAB_1BY5_PACKED_SIZE] = '{
{1'b0,  8'd14,  9'd29},{1'b1,  8'd15, 9'd145},
{1'b0,   8'd3, 9'd172},{1'b1,   8'd7, 9'd255},
{1'b0,   8'd3, 9'd136},{1'b1,   8'd6, 9'd204},
{1'b0,   8'd3, 9'd328},{1'b1,   8'd4, 9'd170},
{1'b0,   8'd5,  9'd59},{1'b1,   8'd8, 9'd287},
{1'b0,   8'd1, 9'd132},{1'b1,   8'd4, 9'd222},
{1'b0,   8'd0, 9'd253},{1'b1,   8'd8, 9'd152},
{1'b0,  8'd10, 9'd304},{1'b1,  8'd16,  9'd10},
{1'b0,   8'd1, 9'd133},{1'b1,   8'd6,   9'd2},
{1'b0,   8'd2, 9'd249},{1'b1,  8'd10,  9'd99},
{1'b0,   8'd2, 9'd158},{1'b1,   8'd9,  9'd95},
{1'b0,   8'd7, 9'd265},{1'b1,  8'd14, 9'd144},
{1'b0,   8'd0,  9'd68},{1'b1,   8'd8, 9'd158},
{1'b0,   8'd4, 9'd307},{1'b1,   8'd8, 9'd335},
{1'b0,   8'd4,  9'd57},{1'b1,   8'd5,  9'd14},
{1'b0,   8'd5, 9'd274},{1'b1,  8'd17, 9'd314},
{1'b0,   8'd1,  9'd85},{1'b1,   8'd4,  9'd58},
{1'b0,   8'd0,  9'd66},{1'b1,   8'd4, 9'd325},
{1'b0,   8'd4, 9'd299},{1'b1,   8'd7, 9'd273},
{1'b0,   8'd0,  9'd93},{1'b1,   8'd6, 9'd230},
{1'b0,   8'd6,  9'd59},{1'b1,   8'd7, 9'd282},
{1'b0,   8'd1,  9'd72},{1'b1,   8'd8, 9'd171},
{1'b0,   8'd1,  9'd28},{1'b1,  8'd12, 9'd228},
{1'b0,   8'd4, 9'd122},{1'b1,   8'd7,  9'd66},
{1'b0,   8'd0, 9'd359},{1'b1,   8'd5, 9'd230},
{1'b0,   8'd3, 9'd220},{1'b1,   8'd5, 9'd257},
{1'b0,   8'd7, 9'd311},{1'b1,   8'd8, 9'd113},
{1'b0,   8'd1,  9'd33},{1'b1,   8'd8, 9'd316},
{1'b0,   8'd8, 9'd273},{1'b1,  8'd13, 9'd208},
{1'b0,   8'd1,   9'd9},{1'b1,   8'd4, 9'd236},
{1'b0,   8'd5,  9'd17},{1'b1,   8'd8, 9'd228},
{1'b0,   8'd0,  9'd62},{1'b1,   8'd7, 9'd152},
{1'b0,   8'd3, 9'd227},{1'b1,   8'd5,  9'd96},
{1'b0,  8'd11, 9'd335},{1'b1,  8'd13, 9'd145},
{1'b0,   8'd9, 9'd236},{1'b1,  8'd15, 9'd186},
{1'b0,   8'd3,  9'd11},{1'b1,   8'd4, 9'd118},
{1'b0,   8'd1, 9'd328},{1'b1,   8'd7,  9'd51},
{1'b0,   8'd5, 9'd247},{1'b1,  8'd12, 9'd109},
{1'b0,   8'd2, 9'd122},{1'b1,   8'd4, 9'd134},
{1'b0,   8'd2, 9'd268},{1'b1,   8'd7,  9'd21},
{1'b0,   8'd0, 9'd299},{1'b1,   8'd2,  9'd61},
{1'b0,   8'd2,   9'd6},{1'b1,   8'd3, 9'd161},
{1'b0,   8'd1, 9'd279},{1'b1,   8'd2, 9'd339},
{1'b0,   8'd3, 9'd262},{1'b1,   8'd5, 9'd273},
{1'b0,   8'd0, 9'd162},{1'b1,   8'd7, 9'd230},
{1'b0,   8'd2, 9'd247},{1'b1,   8'd9,  9'd17},
{1'b0,   8'd2, 9'd202},{1'b1,   8'd6,  9'd98},
{1'b0,   8'd1, 9'd294},{1'b1,   8'd3, 9'd300},
{1'b0,   8'd5,  9'd82},{1'b1,   8'd6, 9'd340},
{1'b0,   8'd6, 9'd359},{1'b1,   8'd7,  9'd80},
{1'b0,   8'd6, 9'd225},{1'b1,  8'd11, 9'd164},
{1'b0,   8'd0, 9'd125},{1'b1,   8'd2,   9'd3},
{1'b0,   8'd2, 9'd306},{1'b1,   8'd6, 9'd326},
{1'b0,   8'd1,  9'd10},{1'b1,   8'd5, 9'd215},
{1'b0,   8'd8, 9'd173},{1'b1,  8'd15, 9'd297},
{1'b0,   8'd7, 9'd101},{1'b1,  8'd11, 9'd184},
{1'b0,  8'd16, 9'd245},{1'b1,  8'd17, 9'd116},
{1'b0,   8'd1, 9'd291},{1'b1,   8'd6,   9'd1},
{1'b0,   8'd1, 9'd289},{1'b1,   8'd3, 9'd171},
{1'b0,   8'd2, 9'd321},{1'b1,  8'd14, 9'd139},
{1'b0,   8'd0, 9'd193},{1'b1,  8'd13, 9'd111},
{1'b0,   8'd6, 9'd137},{1'b1,  8'd12, 9'd177},
{1'b0,   8'd6, 9'd155},{1'b1,   8'd8, 9'd348},
{1'b0,   8'd5, 9'd281},{1'b1,   8'd6,  9'd13},
{1'b0,   8'd0, 9'd264},{1'b1,   8'd2, 9'd276},
{1'b0,   8'd3, 9'd232},{1'b1,  8'd17, 9'd247},
{1'b0,   8'd3, 9'd151},{1'b1,   8'd8, 9'd191},
{1'b0,   8'd0, 9'd308},{1'b1,   8'd5,  9'd43},
{1'b0,   8'd8, 9'd104},{1'b1,  8'd16, 9'd168},
{1'b0,   8'd0, 9'd316},{1'b1,   8'd4, 9'd204},
{1'b0,   8'd7,  9'd47},{1'b1,  8'd10, 9'd350},
{1'b0,   8'd3,  9'd70},{1'b1,   8'd4, 9'd105}
};
localparam int          cMEDIUM_HS_TAB_11BY45_PACKED_SIZE = 136;
localparam bit [17 : 0] cMEDIUM_HS_TAB_11BY45_PACKED[cMEDIUM_HS_TAB_11BY45_PACKED_SIZE] = '{
{1'b0,  8'd10,  9'd67},{1'b1,  8'd21,  9'd58},
{1'b0,   8'd2, 9'd158},{1'b1,   8'd7, 9'd296},
{1'b0,  8'd15, 9'd168},{1'b1,  8'd17, 9'd262},
{1'b0,   8'd0, 9'd253},{1'b1,   8'd3, 9'd140},
{1'b0,   8'd8,  9'd85},{1'b1,   8'd9, 9'd259},
{1'b0,   8'd1, 9'd248},{1'b1,   8'd5,  9'd21},
{1'b0,   8'd0, 9'd176},{1'b1,   8'd7, 9'd177},
{1'b0,   8'd7, 9'd173},{1'b1,  8'd21, 9'd192},
{1'b0,   8'd3, 9'd206},{1'b1,   8'd5,  9'd32},
{1'b0,   8'd3, 9'd241},{1'b1,   8'd4,  9'd66},
{1'b0,   8'd2, 9'd209},{1'b1,  8'd11, 9'd172},
{1'b0,  8'd13,  9'd39},{1'b1,  8'd20, 9'd156},
{1'b0,  8'd16,  9'd78},{1'b1,  8'd21,  9'd83},
{1'b0,   8'd0, 9'd303},{1'b1,   8'd5,  9'd57},
{1'b0,   8'd9, 9'd248},{1'b1,  8'd15, 9'd291},
{1'b0,   8'd1, 9'd197},{1'b1,   8'd4, 9'd277},
{1'b0,   8'd4, 9'd211},{1'b1,   8'd5, 9'd256},
{1'b0,   8'd3, 9'd275},{1'b1,   8'd6,   9'd6},
{1'b0,   8'd2,  9'd34},{1'b1,   8'd8, 9'd129},
{1'b0,   8'd9, 9'd234},{1'b1,  8'd12,  9'd37},
{1'b0,   8'd9,  9'd85},{1'b1,  8'd14, 9'd103},
{1'b0,   8'd0, 9'd218},{1'b1,   8'd8, 9'd260},
{1'b0,   8'd1, 9'd218},{1'b1,   8'd5, 9'd314},
{1'b0,   8'd6,  9'd30},{1'b1,  8'd10, 9'd320},
{1'b0,   8'd2, 9'd347},{1'b1,   8'd7, 9'd341},
{1'b0,   8'd7, 9'd141},{1'b1,  8'd16, 9'd181},
{1'b0,   8'd6, 9'd329},{1'b1,  8'd12, 9'd228},
{1'b0,   8'd0, 9'd235},{1'b1,   8'd1,  9'd37},
{1'b0,   8'd1, 9'd315},{1'b1,  8'd10,  9'd22},
{1'b0,   8'd3, 9'd139},{1'b1,  8'd17, 9'd169},
{1'b0,   8'd5,  9'd20},{1'b1,  8'd16, 9'd234},
{1'b0,   8'd6, 9'd307},{1'b1,   8'd8, 9'd307},
{1'b0,   8'd2,  9'd76},{1'b1,   8'd3, 9'd320},
{1'b0,   8'd1, 9'd299},{1'b1,   8'd2,  9'd95},
{1'b0,   8'd6, 9'd217},{1'b1,   8'd7, 9'd314},
{1'b0,   8'd4,  9'd94},{1'b1,   8'd9, 9'd104},
{1'b0,   8'd4,  9'd60},{1'b1,   8'd5, 9'd258},
{1'b0,   8'd6,  9'd65},{1'b1,  8'd19, 9'd191},
{1'b0,   8'd8, 9'd316},{1'b1,   8'd9, 9'd289},
{1'b0,   8'd2, 9'd303},{1'b1,   8'd7, 9'd122},
{1'b0,   8'd0,  9'd59},{1'b1,  8'd11, 9'd295},
{1'b0,   8'd1, 9'd244},{1'b1,   8'd4,  9'd55},
{1'b0,  8'd13, 9'd177},{1'b1,  8'd17,  9'd46},
{1'b0,   8'd6,  9'd10},{1'b1,   8'd8, 9'd218},
{1'b0,   8'd5, 9'd188},{1'b1,   8'd6, 9'd103},
{1'b0,  8'd14, 9'd288},{1'b1,  8'd18,  9'd33},
{1'b0,   8'd4, 9'd259},{1'b1,   8'd9,  9'd11},
{1'b0,   8'd1,  9'd11},{1'b1,   8'd5, 9'd152},
{1'b0,   8'd8, 9'd282},{1'b1,  8'd18, 9'd349},
{1'b0,   8'd7, 9'd239},{1'b1,   8'd9, 9'd139},
{1'b0,  8'd14, 9'd297},{1'b1,  8'd20, 9'd150},
{1'b0,   8'd8, 9'd260},{1'b1,  8'd18, 9'd243},
{1'b0,   8'd7, 9'd141},{1'b1,  8'd15, 9'd172},
{1'b0,   8'd3, 9'd187},{1'b1,  8'd19,  9'd97},
{1'b0,   8'd0,   9'd2},{1'b1,   8'd2, 9'd216},
{1'b0,   8'd0, 9'd331},{1'b1,   8'd2,  9'd40},
{1'b0,   8'd1, 9'd343},{1'b1,   8'd3, 9'd107},
{1'b0,   8'd7, 9'd198},{1'b1,   8'd8, 9'd183},
{1'b0,   8'd4, 9'd337},{1'b1,  8'd20, 9'd294},
{1'b0,  8'd13,  9'd56},{1'b1,  8'd19, 9'd249},
{1'b0,   8'd5, 9'd307},{1'b1,   8'd6,  9'd59},
{1'b0,   8'd3, 9'd138},{1'b1,   8'd6, 9'd138},
{1'b0,   8'd0, 9'd108},{1'b1,   8'd3, 9'd325},
{1'b0,   8'd2, 9'd307},{1'b1,   8'd9, 9'd257},
{1'b0,   8'd9, 9'd342},{1'b1,  8'd12,  9'd89},
{1'b0,   8'd1, 9'd291},{1'b1,   8'd4,  9'd37},
{1'b0,   8'd4,  9'd42},{1'b1,   8'd8,  9'd15},
{1'b0,   8'd0, 9'd100},{1'b1,  8'd11, 9'd347}
};
localparam int          cMEDIUM_HS_TAB_1BY3_PACKED_SIZE = 180;
localparam bit [17 : 0] cMEDIUM_HS_TAB_1BY3_PACKED[cMEDIUM_HS_TAB_1BY3_PACKED_SIZE] = '{
{1'b0,   8'd1, 9'd219},{1'b0,   8'd2, 9'd256},{1'b1,   8'd3, 9'd212},
{1'b0,   8'd3,  9'd69},{1'b0,   8'd8, 9'd144},{1'b1,  8'd23,  9'd83},
{1'b0,   8'd4, 9'd253},{1'b0,   8'd7, 9'd234},{1'b1,   8'd9, 9'd226},
{1'b0,   8'd0,  9'd17},{1'b0,   8'd5, 9'd296},{1'b1,  8'd11,  9'd62},
{1'b0,   8'd5,  9'd86},{1'b0,  8'd24, 9'd356},{1'b1,  8'd28,  9'd37},
{1'b0,   8'd7, 9'd100},{1'b0,  8'd18, 9'd134},{1'b1,  8'd21, 9'd265},
{1'b0,   8'd0, 9'd343},{1'b0,  8'd23, 9'd269},{1'b1,  8'd26, 9'd104},
{1'b0,   8'd8,  9'd50},{1'b0,   8'd9,  9'd14},{1'b1,  8'd10, 9'd313},
{1'b0,   8'd7,  9'd56},{1'b0,   8'd8, 9'd136},{1'b1,  8'd17, 9'd110},
{1'b0,   8'd2,  9'd55},{1'b0,   8'd5, 9'd320},{1'b1,   8'd6, 9'd143},
{1'b0,   8'd1,  9'd35},{1'b0,   8'd9,  9'd92},{1'b1,  8'd14, 9'd233},
{1'b0,   8'd4,  9'd94},{1'b0,  8'd22, 9'd129},{1'b1,  8'd25,  9'd34},
{1'b0,   8'd4, 9'd338},{1'b0,   8'd5, 9'd232},{1'b1,  8'd15, 9'd173},
{1'b0,   8'd0,  9'd68},{1'b0,   8'd7, 9'd267},{1'b1,   8'd8,  9'd48},
{1'b0,   8'd3,  9'd58},{1'b0,   8'd6, 9'd272},{1'b1,  8'd16, 9'd317},
{1'b0,   8'd6,  9'd12},{1'b0,   8'd9, 9'd245},{1'b1,  8'd14, 9'd114},
{1'b0,   8'd2,  9'd53},{1'b0,   8'd8,  9'd26},{1'b1,  8'd22, 9'd275},
{1'b0,   8'd1,  9'd54},{1'b0,   8'd2,  9'd46},{1'b1,   8'd5,  9'd21},
{1'b0,   8'd1, 9'd250},{1'b0,   8'd5,  9'd20},{1'b1,   8'd7,  9'd96},
{1'b0,   8'd7,  9'd11},{1'b0,  8'd18, 9'd328},{1'b1,  8'd19, 9'd120},
{1'b0,   8'd3,  9'd23},{1'b0,   8'd4,  9'd64},{1'b1,   8'd9, 9'd312},
{1'b0,   8'd3, 9'd303},{1'b0,   8'd6, 9'd228},{1'b1,   8'd9, 9'd164},
{1'b0,   8'd6,  9'd91},{1'b0,   8'd8, 9'd275},{1'b1,  8'd11,  9'd40},
{1'b0,   8'd1,  9'd50},{1'b0,   8'd2, 9'd100},{1'b1,   8'd4,  9'd32},
{1'b0,   8'd0, 9'd271},{1'b0,   8'd5,  9'd95},{1'b1,  8'd13,  9'd51},
{1'b0,   8'd0, 9'd292},{1'b0,   8'd5, 9'd298},{1'b1,   8'd8, 9'd175},
{1'b0,   8'd2, 9'd239},{1'b0,  8'd12, 9'd223},{1'b1,  8'd20, 9'd329},
{1'b0,   8'd3, 9'd137},{1'b0,   8'd6,  9'd94},{1'b1,  8'd10, 9'd174},
{1'b0,   8'd1, 9'd231},{1'b0,   8'd4, 9'd115},{1'b1,   8'd9, 9'd290},
{1'b0,   8'd7, 9'd297},{1'b0,  8'd11, 9'd179},{1'b1,  8'd13,  9'd99},
{1'b0,   8'd6,  9'd82},{1'b0,   8'd8, 9'd184},{1'b1,  8'd23, 9'd337},
{1'b0,   8'd1, 9'd315},{1'b0,   8'd2, 9'd111},{1'b1,  8'd15, 9'd172},
{1'b0,   8'd2,  9'd73},{1'b0,   8'd5,  9'd98},{1'b1,  8'd27, 9'd277},
{1'b0,   8'd0, 9'd168},{1'b0,   8'd4,  9'd44},{1'b1,   8'd9, 9'd186},
{1'b0,   8'd3, 9'd188},{1'b0,  8'd22, 9'd142},{1'b1,  8'd28,  9'd94},
{1'b0,   8'd3,  9'd52},{1'b0,   8'd5, 9'd342},{1'b1,  8'd12, 9'd133},
{1'b0,   8'd0, 9'd123},{1'b0,   8'd7,  9'd45},{1'b1,  8'd10, 9'd102},
{1'b0,   8'd1,  9'd25},{1'b0,   8'd8,  9'd11},{1'b1,  8'd29, 9'd187},
{1'b0,   8'd1,  9'd26},{1'b0,   8'd4, 9'd350},{1'b1,  8'd19,  9'd76},
{1'b0,   8'd0, 9'd203},{1'b0,   8'd2,   9'd5},{1'b1,   8'd4, 9'd215},
{1'b0,   8'd2, 9'd289},{1'b0,   8'd5, 9'd103},{1'b1,   8'd9, 9'd169},
{1'b0,   8'd7, 9'd169},{1'b0,  8'd21, 9'd293},{1'b1,  8'd26, 9'd128},
{1'b0,   8'd0, 9'd278},{1'b0,  8'd25, 9'd147},{1'b1,  8'd27,  9'd91},
{1'b0,   8'd8, 9'd238},{1'b0,  8'd25, 9'd284},{1'b1,  8'd27, 9'd300},
{1'b0,   8'd6, 9'd205},{1'b0,  8'd14,  9'd62},{1'b1,  8'd24, 9'd208},
{1'b0,   8'd1, 9'd231},{1'b0,   8'd3,  9'd47},{1'b1,   8'd6, 9'd110},
{1'b0,   8'd4, 9'd108},{1'b0,   8'd7, 9'd291},{1'b1,   8'd8, 9'd128},
{1'b0,   8'd7, 9'd296},{1'b0,  8'd17, 9'd195},{1'b1,  8'd21, 9'd124},
{1'b0,   8'd3, 9'd198},{1'b0,  8'd17,  9'd69},{1'b1,  8'd18, 9'd148},
{1'b0,   8'd0, 9'd330},{1'b0,   8'd9,  9'd82},{1'b1,  8'd13, 9'd265},
{1'b0,   8'd2, 9'd117},{1'b0,   8'd6, 9'd319},{1'b1,   8'd9, 9'd287},
{1'b0,   8'd6, 9'd253},{1'b0,  8'd19, 9'd189},{1'b1,  8'd20, 9'd197},
{1'b0,  8'd20,  9'd94},{1'b0,  8'd28,  9'd23},{1'b1,  8'd29,  9'd21},
{1'b0,   8'd5, 9'd103},{1'b0,  8'd24, 9'd179},{1'b1,  8'd29, 9'd140},
{1'b0,   8'd0,  9'd25},{1'b0,   8'd1,  9'd16},{1'b1,   8'd3, 9'd293},
{1'b0,   8'd0, 9'd152},{1'b0,   8'd7, 9'd137},{1'b1,  8'd26,  9'd21},
{1'b0,   8'd4,   9'd5},{1'b0,   8'd9, 9'd321},{1'b1,  8'd12, 9'd311},
{1'b0,   8'd1, 9'd176},{1'b0,   8'd3, 9'd267},{1'b1,   8'd4,  9'd65},
{1'b0,   8'd2, 9'd305},{1'b0,   8'd6,  9'd74},{1'b1,  8'd16, 9'd267},
{1'b0,   8'd8, 9'd170},{1'b0,  8'd15, 9'd262},{1'b1,  8'd16, 9'd187}
};
