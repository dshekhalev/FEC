//
// Project       : polar code 3gpp
// Author        : Shekhalev Denis (des00)
// Workfile      : pc_3ggp_ts_38_212_tab.svh
// Description   : Reliability table for bit channel from 3GPP TS 38.212 V15.1.1 (2018-4)
//

localparam int bits_addr_tab [1024] = '{1023, 1022, 1021, 1019, 1015, 1007, 1020, 991, 1018, 1017, 1014, 1006, 895, 1013, 1011, 959, 1005, 990, 1003, 989, 767, 1016, 999, 1012, 987, 958, 983, 957, 1010, 1004, 955, 1009, 894, 975, 893, 1002, 951, 1001, 988, 511, 766, 998, 891, 943, 986, 997, 985, 887, 956, 765, 995, 927, 982, 981, 879, 954, 974, 763, 953, 979, 510, 1008, 759, 863, 950, 892, 1000, 973, 949, 509, 890, 971, 996, 942, 751, 984, 889, 507, 947, 831, 886, 967, 941, 764, 926, 980, 994, 939, 885, 993, 735, 878, 925, 503, 762, 883, 978, 935, 703, 495, 952, 877, 761, 972, 923, 977, 948, 758, 862, 875, 919, 970, 757, 861, 508, 969, 750, 946, 479, 888, 639, 871, 911, 830, 940, 859, 755, 966, 945, 749, 506, 884, 938, 965, 829, 734, 924, 855, 505, 747, 963, 937, 882, 934, 827, 733, 447, 992, 847, 876, 501, 921, 702, 494, 881, 760, 743, 933, 502, 918, 874, 922, 823, 731, 499, 860, 756, 931, 701, 873, 493, 727, 917, 870, 976, 815, 910, 383, 968, 478, 858, 754, 699, 491, 869, 944, 748, 638, 915, 477, 719, 909, 964, 255, 799, 504, 857, 854, 753, 828, 746, 695, 487, 907, 637, 867, 853, 475, 936, 962, 446, 732, 826, 745, 846, 500, 825, 903, 687, 932, 635, 471, 445, 742, 880, 498, 730, 851, 822, 382, 920, 845, 741, 443, 700, 729, 631, 492, 872, 961, 726, 821, 930, 497, 381, 843, 463, 916, 739, 671, 623, 490, 929, 439, 814, 819, 868, 752, 914, 698, 725, 839, 856, 476, 813, 718, 908, 486, 723, 866, 489, 607, 431, 697, 379, 811, 798, 913, 575, 717, 254, 694, 636, 474, 807, 715, 906, 797, 693, 865, 960, 852, 744, 634, 473, 795, 905, 485, 415, 483, 470, 444, 375, 850, 740, 686, 902, 824, 691, 253, 711, 633, 844, 685, 630, 901, 367, 791, 928, 728, 820, 849, 783, 670, 899, 738, 842, 683, 247, 469, 441, 442, 462, 251, 737, 438, 467, 351, 629, 841, 724, 679, 669, 496, 461, 818, 380, 437, 627, 622, 459, 378, 239, 488, 667, 838, 430, 484, 812, 621, 319, 817, 435, 377, 696, 722, 912, 606, 810, 864, 716, 837, 721, 714, 809, 796, 455, 472, 619, 835, 692, 663, 223, 414, 904, 427, 806, 482, 632, 713, 690, 848, 605, 373, 252, 794, 429, 710, 684, 615, 805, 900, 655, 468, 366, 603, 413, 574, 481, 371, 250, 793, 466, 423, 374, 689, 628, 440, 365, 709, 789, 803, 411, 573, 682, 249, 460, 790, 668, 599, 350, 707, 246, 681, 465, 571, 626, 436, 407, 782, 191, 127, 363, 620, 666, 458, 245, 349, 677, 434, 678, 591, 787, 399, 457, 359, 238, 625, 840, 567, 736, 665, 428, 376, 781, 898, 618, 675, 318, 454, 662, 243, 897, 347, 836, 816, 720, 433, 604, 617, 779, 808, 661, 834, 712, 804, 833, 559, 237, 453, 426, 222, 317, 775, 372, 343, 412, 235, 543, 614, 451, 425, 422, 613, 370, 221, 315, 480, 335, 659, 654, 364, 190, 369, 248, 653, 688, 231, 410, 602, 611, 802, 792, 421, 651, 601, 598, 708, 311, 219, 572, 597, 788, 570, 409, 590, 362, 801, 680, 464, 406, 419, 348, 647, 786, 215, 589, 706, 361, 676, 566, 189, 595, 244, 569, 303, 405, 358, 456, 346, 398, 565, 242, 126, 705, 780, 587, 624, 664, 236, 187, 357, 432, 785, 558, 674, 207, 403, 397, 452, 345, 563, 778, 241, 316, 342, 616, 660, 557, 125, 234, 183, 287, 355, 583, 673, 395, 424, 314, 220, 777, 341, 612, 658, 123, 175, 774, 555, 233, 334, 542, 450, 313, 391, 230, 652, 368, 218, 339, 600, 119, 333, 657, 610, 773, 541, 310, 420, 159, 229, 650, 551, 596, 609, 408, 217, 449, 188, 309, 214, 331, 111, 539, 360, 771, 649, 302, 418, 594, 896, 227, 404, 646, 186, 588, 832, 568, 213, 417, 301, 307, 356, 402, 800, 564, 327, 95, 206, 240, 535, 593, 645, 586, 344, 396, 185, 401, 211, 354, 299, 585, 286, 562, 643, 182, 205, 124, 232, 285, 295, 181, 556, 582, 527, 394, 340, 63, 203, 561, 353, 448, 122, 283, 393, 581, 554, 174, 390, 704, 312, 338, 228, 179, 784, 199, 553, 121, 173, 389, 540, 579, 332, 118, 672, 550, 337, 158, 279, 271, 416, 216, 308, 387, 538, 549, 226, 330, 776, 171, 212, 117, 110, 329, 656, 157, 772, 306, 326, 225, 167, 115, 537, 534, 184, 109, 300, 547, 305, 210, 155, 533, 325, 352, 608, 400, 298, 204, 94, 648, 284, 209, 151, 180, 107, 770, 297, 392, 323, 592, 202, 644, 93, 294, 178, 103, 143, 282, 62, 336, 201, 120, 172, 198, 769, 584, 91, 388, 293, 177, 526, 278, 281, 642, 525, 531, 61, 170, 116, 197, 87, 156, 277, 114, 560, 169, 59, 291, 580, 275, 523, 641, 270, 195, 552, 519, 166, 224, 578, 108, 269, 79, 154, 113, 548, 577, 536, 328, 55, 106, 165, 153, 150, 386, 208, 324, 546, 385, 267, 47, 92, 163, 296, 304, 105, 102, 149, 263, 532, 322, 292, 545, 90, 200, 31, 321, 530, 142, 176, 147, 101, 141, 196, 524, 529, 290, 89, 280, 60, 86, 99, 139, 168, 58, 522, 276, 85, 194, 289, 78, 135, 112, 521, 57, 83, 54, 518, 274, 268, 768, 164, 77, 152, 193, 53, 162, 104, 517, 273, 266, 75, 46, 148, 51, 640, 100, 45, 576, 161, 265, 262, 71, 146, 30, 140, 88, 515, 98, 43, 29, 261, 145, 138, 84, 259, 39, 97, 27, 56, 82, 137, 76, 384, 134, 23, 52, 133, 320, 15, 73, 50, 81, 131, 44, 70, 544, 192, 528, 288, 520, 160, 272, 74, 49, 516, 42, 69, 28, 144, 41, 67, 96, 514, 38, 264, 260, 136, 22, 25, 37, 80, 513, 26, 258, 35, 132, 21, 257, 72, 14, 48, 13, 19, 130, 68, 40, 11, 512, 66, 129, 7, 36, 24, 34, 256, 20, 65, 33, 12, 128, 18, 10, 17, 6, 9, 64, 5, 3, 32, 16, 8, 4, 2, 1, 0};
