//
// (!!!) IT'S GENERATED short table for 7/8 coderate, 8176 bits do 7 LLR per cycle(!!!)
//
  addr_tab[0][0][0][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6}, invsela:'{0, 1, 2, 3, 4, 5, 6}};
  addr_tab[0][0][1][0] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 2047, 2047}, offsetm:'{0, 0, 0, 0, 0, 2047, 2047}, sela:'{5, 6, 0, 1, 2, 3, 4}, invsela:'{2, 3, 4, 5, 6, 0, 1}};
  addr_tab[0][0][2][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6}, invsela:'{0, 1, 2, 3, 4, 5, 6}};
  addr_tab[0][0][3][0] = '{baddr:4, offset:'{0, 0, 0, 2047, 2047, 2047, 2047}, offsetm:'{0, 0, 0, 2047, 2047, 2047, 2047}, sela:'{3, 4, 5, 6, 0, 1, 2}, invsela:'{4, 5, 6, 0, 1, 2, 3}};
  addr_tab[0][0][4][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6}, invsela:'{0, 1, 2, 3, 4, 5, 6}};
  addr_tab[0][0][5][0] = '{baddr:22, offset:'{0, 0, 0, 0, 2047, 2047, 2047}, offsetm:'{0, 0, 0, 0, 2047, 2047, 2047}, sela:'{4, 5, 6, 0, 1, 2, 3}, invsela:'{3, 4, 5, 6, 0, 1, 2}};
  addr_tab[0][0][6][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6}, invsela:'{0, 1, 2, 3, 4, 5, 6}};
  addr_tab[0][0][7][0] = '{baddr:2, offset:'{0, 0, 2047, 2047, 2047, 2047, 2047}, offsetm:'{0, 0, 2047, 2047, 2047, 2047, 2047}, sela:'{2, 3, 4, 5, 6, 0, 1}, invsela:'{5, 6, 0, 1, 2, 3, 4}};
  addr_tab[0][0][8][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6}, invsela:'{0, 1, 2, 3, 4, 5, 6}};
  addr_tab[0][0][9][0] = '{baddr:8, offset:'{0, 0, 0, 0, 2047, 2047, 2047}, offsetm:'{0, 0, 0, 0, 2047, 2047, 2047}, sela:'{4, 5, 6, 0, 1, 2, 3}, invsela:'{3, 4, 5, 6, 0, 1, 2}};
  addr_tab[0][0][10][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6}, invsela:'{0, 1, 2, 3, 4, 5, 6}};
  addr_tab[0][0][11][0] = '{baddr:3, offset:'{0, 0, 0, 0, 2047, 2047, 2047}, offsetm:'{0, 0, 0, 0, 2047, 2047, 2047}, sela:'{4, 5, 6, 0, 1, 2, 3}, invsela:'{3, 4, 5, 6, 0, 1, 2}};
  addr_tab[0][0][12][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6}, invsela:'{0, 1, 2, 3, 4, 5, 6}};
  addr_tab[0][0][13][0] = '{baddr:29, offset:'{0, 0, 0, 0, 0, 0, 2047}, offsetm:'{0, 0, 0, 0, 0, 0, 2047}, sela:'{6, 0, 1, 2, 3, 4, 5}, invsela:'{1, 2, 3, 4, 5, 6, 0}};
  addr_tab[0][0][14][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6}, invsela:'{0, 1, 2, 3, 4, 5, 6}};
  addr_tab[0][0][15][0] = '{baddr:6, offset:'{0, 2047, 2047, 2047, 2047, 2047, 2047}, offsetm:'{0, 2047, 2047, 2047, 2047, 2047, 2047}, sela:'{1, 2, 3, 4, 5, 6, 0}, invsela:'{6, 0, 1, 2, 3, 4, 5}};
  addr_tab[0][1][0][0] = '{baddr:26, offset:'{0, 2047, 2047, 2047, 2047, 2047, 2047}, offsetm:'{0, 2047, 2047, 2047, 2047, 2047, 2047}, sela:'{1, 2, 3, 4, 5, 6, 0}, invsela:'{6, 0, 1, 2, 3, 4, 5}};
  addr_tab[0][1][1][0] = '{baddr:35, offset:'{0, 2047, 2047, 2047, 2047, 2047, 2047}, offsetm:'{0, 2047, 2047, 2047, 2047, 2047, 2047}, sela:'{1, 2, 3, 4, 5, 6, 0}, invsela:'{6, 0, 1, 2, 3, 4, 5}};
  addr_tab[0][1][2][0] = '{baddr:51, offset:'{0, 0, 2047, 2047, 2047, 2047, 2047}, offsetm:'{0, 0, 2047, 2047, 2047, 2047, 2047}, sela:'{2, 3, 4, 5, 6, 0, 1}, invsela:'{5, 6, 0, 1, 2, 3, 4}};
  addr_tab[0][1][3][0] = '{baddr:62, offset:'{0, 0, 0, 0, 2047, 2047, 2047}, offsetm:'{0, 0, 0, 0, 2047, 2047, 2047}, sela:'{4, 5, 6, 0, 1, 2, 3}, invsela:'{3, 4, 5, 6, 0, 1, 2}};
  addr_tab[0][1][4][0] = '{baddr:56, offset:'{0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6}, invsela:'{0, 1, 2, 3, 4, 5, 6}};
  addr_tab[0][1][5][0] = '{baddr:59, offset:'{0, 0, 0, 2047, 2047, 2047, 2047}, offsetm:'{0, 0, 0, 2047, 2047, 2047, 2047}, sela:'{3, 4, 5, 6, 0, 1, 2}, invsela:'{4, 5, 6, 0, 1, 2, 3}};
  addr_tab[0][1][6][0] = '{baddr:51, offset:'{0, 2047, 2047, 2047, 2047, 2047, 2047}, offsetm:'{0, 2047, 2047, 2047, 2047, 2047, 2047}, sela:'{1, 2, 3, 4, 5, 6, 0}, invsela:'{6, 0, 1, 2, 3, 4, 5}};
  addr_tab[0][1][7][0] = '{baddr:52, offset:'{0, 0, 2047, 2047, 2047, 2047, 2047}, offsetm:'{0, 0, 2047, 2047, 2047, 2047, 2047}, sela:'{2, 3, 4, 5, 6, 0, 1}, invsela:'{5, 6, 0, 1, 2, 3, 4}};
  addr_tab[0][1][8][0] = '{baddr:44, offset:'{0, 0, 0, 0, 0, 0, 2047}, offsetm:'{0, 0, 0, 0, 0, 0, 2047}, sela:'{6, 0, 1, 2, 3, 4, 5}, invsela:'{1, 2, 3, 4, 5, 6, 0}};
  addr_tab[0][1][9][0] = '{baddr:47, offset:'{0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6}, invsela:'{0, 1, 2, 3, 4, 5, 6}};
  addr_tab[0][1][10][0] = '{baddr:30, offset:'{0, 0, 0, 0, 2047, 2047, 2047}, offsetm:'{0, 0, 0, 0, 2047, 2047, 2047}, sela:'{4, 5, 6, 0, 1, 2, 3}, invsela:'{3, 4, 5, 6, 0, 1, 2}};
  addr_tab[0][1][11][0] = '{baddr:41, offset:'{0, 2047, 2047, 2047, 2047, 2047, 2047}, offsetm:'{0, 2047, 2047, 2047, 2047, 2047, 2047}, sela:'{1, 2, 3, 4, 5, 6, 0}, invsela:'{6, 0, 1, 2, 3, 4, 5}};
  addr_tab[0][1][12][0] = '{baddr:57, offset:'{0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6}, invsela:'{0, 1, 2, 3, 4, 5, 6}};
  addr_tab[0][1][13][0] = '{baddr:66, offset:'{0, 0, 2047, 2047, 2047, 2047, 2047}, offsetm:'{0, 0, 2047, 2047, 2047, 2047, 2047}, sela:'{2, 3, 4, 5, 6, 0, 1}, invsela:'{5, 6, 0, 1, 2, 3, 4}};
  addr_tab[0][1][14][0] = '{baddr:36, offset:'{0, 0, 2047, 2047, 2047, 2047, 2047}, offsetm:'{0, 0, 2047, 2047, 2047, 2047, 2047}, sela:'{2, 3, 4, 5, 6, 0, 1}, invsela:'{5, 6, 0, 1, 2, 3, 4}};
  addr_tab[0][1][15][0] = '{baddr:38, offset:'{0, 0, 2047, 2047, 2047, 2047, 2047}, offsetm:'{0, 0, 2047, 2047, 2047, 2047, 2047}, sela:'{2, 3, 4, 5, 6, 0, 1}, invsela:'{5, 6, 0, 1, 2, 3, 4}};
  addr_tab[1][0][0][0] = '{baddr:15, offset:'{0, 2047, 2047, 2047, 2047, 2047, 2047}, offsetm:'{0, 2047, 2047, 2047, 2047, 2047, 2047}, sela:'{1, 2, 3, 4, 5, 6, 0}, invsela:'{6, 0, 1, 2, 3, 4, 5}};
  addr_tab[1][0][1][0] = '{baddr:19, offset:'{0, 0, 0, 0, 2047, 2047, 2047}, offsetm:'{0, 0, 0, 0, 2047, 2047, 2047}, sela:'{4, 5, 6, 0, 1, 2, 3}, invsela:'{3, 4, 5, 6, 0, 1, 2}};
  addr_tab[1][0][2][0] = '{baddr:29, offset:'{0, 0, 2047, 2047, 2047, 2047, 2047}, offsetm:'{0, 0, 2047, 2047, 2047, 2047, 2047}, sela:'{2, 3, 4, 5, 6, 0, 1}, invsela:'{5, 6, 0, 1, 2, 3, 4}};
  addr_tab[1][0][3][0] = '{baddr:38, offset:'{0, 2047, 2047, 2047, 2047, 2047, 2047}, offsetm:'{0, 2047, 2047, 2047, 2047, 2047, 2047}, sela:'{1, 2, 3, 4, 5, 6, 0}, invsela:'{6, 0, 1, 2, 3, 4, 5}};
  addr_tab[1][0][4][0] = '{baddr:31, offset:'{0, 0, 0, 0, 0, 2047, 2047}, offsetm:'{0, 0, 0, 0, 0, 2047, 2047}, sela:'{5, 6, 0, 1, 2, 3, 4}, invsela:'{2, 3, 4, 5, 6, 0, 1}};
  addr_tab[1][0][5][0] = '{baddr:41, offset:'{0, 0, 2047, 2047, 2047, 2047, 2047}, offsetm:'{0, 0, 2047, 2047, 2047, 2047, 2047}, sela:'{2, 3, 4, 5, 6, 0, 1}, invsela:'{5, 6, 0, 1, 2, 3, 4}};
  addr_tab[1][0][6][0] = '{baddr:7, offset:'{0, 0, 0, 0, 0, 0, 2047}, offsetm:'{0, 0, 0, 0, 0, 0, 2047}, sela:'{6, 0, 1, 2, 3, 4, 5}, invsela:'{1, 2, 3, 4, 5, 6, 0}};
  addr_tab[1][0][7][0] = '{baddr:28, offset:'{0, 0, 0, 0, 2047, 2047, 2047}, offsetm:'{0, 0, 0, 0, 2047, 2047, 2047}, sela:'{4, 5, 6, 0, 1, 2, 3}, invsela:'{3, 4, 5, 6, 0, 1, 2}};
  addr_tab[1][0][8][0] = '{baddr:39, offset:'{0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6}, invsela:'{0, 1, 2, 3, 4, 5, 6}};
  addr_tab[1][0][9][0] = '{baddr:44, offset:'{0, 2047, 2047, 2047, 2047, 2047, 2047}, offsetm:'{0, 2047, 2047, 2047, 2047, 2047, 2047}, sela:'{1, 2, 3, 4, 5, 6, 0}, invsela:'{6, 0, 1, 2, 3, 4, 5}};
  addr_tab[1][0][10][0] = '{baddr:14, offset:'{0, 0, 0, 0, 0, 2047, 2047}, offsetm:'{0, 0, 0, 0, 0, 2047, 2047}, sela:'{5, 6, 0, 1, 2, 3, 4}, invsela:'{2, 3, 4, 5, 6, 0, 1}};
  addr_tab[1][0][11][0] = '{baddr:28, offset:'{0, 0, 2047, 2047, 2047, 2047, 2047}, offsetm:'{0, 0, 2047, 2047, 2047, 2047, 2047}, sela:'{2, 3, 4, 5, 6, 0, 1}, invsela:'{5, 6, 0, 1, 2, 3, 4}};
  addr_tab[1][0][12][0] = '{baddr:35, offset:'{0, 0, 0, 0, 0, 0, 2047}, offsetm:'{0, 0, 0, 0, 0, 0, 2047}, sela:'{6, 0, 1, 2, 3, 4, 5}, invsela:'{1, 2, 3, 4, 5, 6, 0}};
  addr_tab[1][0][13][0] = '{baddr:52, offset:'{0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6}, invsela:'{0, 1, 2, 3, 4, 5, 6}};
  addr_tab[1][0][14][0] = '{baddr:8, offset:'{0, 0, 2047, 2047, 2047, 2047, 2047}, offsetm:'{0, 0, 2047, 2047, 2047, 2047, 2047}, sela:'{2, 3, 4, 5, 6, 0, 1}, invsela:'{5, 6, 0, 1, 2, 3, 4}};
  addr_tab[1][0][15][0] = '{baddr:28, offset:'{0, 0, 0, 2047, 2047, 2047, 2047}, offsetm:'{0, 0, 0, 2047, 2047, 2047, 2047}, sela:'{3, 4, 5, 6, 0, 1, 2}, invsela:'{4, 5, 6, 0, 1, 2, 3}};
  addr_tab[1][1][0][0] = '{baddr:68, offset:'{0, 0, 2047, 2047, 2047, 2047, 2047}, offsetm:'{0, 0, 2047, 2047, 2047, 2047, 2047}, sela:'{2, 3, 4, 5, 6, 0, 1}, invsela:'{5, 6, 0, 1, 2, 3, 4}};
  addr_tab[1][1][1][0] = '{baddr:68, offset:'{0, 0, 0, 0, 2047, 2047, 2047}, offsetm:'{0, 0, 0, 0, 2047, 2047, 2047}, sela:'{4, 5, 6, 0, 1, 2, 3}, invsela:'{3, 4, 5, 6, 0, 1, 2}};
  addr_tab[1][1][2][0] = '{baddr:63, offset:'{0, 2047, 2047, 2047, 2047, 2047, 2047}, offsetm:'{0, 2047, 2047, 2047, 2047, 2047, 2047}, sela:'{1, 2, 3, 4, 5, 6, 0}, invsela:'{6, 0, 1, 2, 3, 4, 5}};
  addr_tab[1][1][3][0] = '{baddr:69, offset:'{0, 0, 2047, 2047, 2047, 2047, 2047}, offsetm:'{0, 0, 2047, 2047, 2047, 2047, 2047}, sela:'{2, 3, 4, 5, 6, 0, 1}, invsela:'{5, 6, 0, 1, 2, 3, 4}};
  addr_tab[1][1][4][0] = '{baddr:60, offset:'{0, 0, 0, 0, 0, 0, 0}, offsetm:'{0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6}, invsela:'{0, 1, 2, 3, 4, 5, 6}};
  addr_tab[1][1][5][0] = '{baddr:69, offset:'{0, 0, 0, 0, 0, 2047, 2047}, offsetm:'{0, 0, 0, 0, 0, 2047, 2047}, sela:'{5, 6, 0, 1, 2, 3, 4}, invsela:'{2, 3, 4, 5, 6, 0, 1}};
  addr_tab[1][1][6][0] = '{baddr:57, offset:'{0, 0, 0, 0, 2047, 2047, 2047}, offsetm:'{0, 0, 0, 0, 2047, 2047, 2047}, sela:'{4, 5, 6, 0, 1, 2, 3}, invsela:'{3, 4, 5, 6, 0, 1, 2}};
  addr_tab[1][1][7][0] = '{baddr:64, offset:'{0, 0, 0, 0, 2047, 2047, 2047}, offsetm:'{0, 0, 0, 0, 2047, 2047, 2047}, sela:'{4, 5, 6, 0, 1, 2, 3}, invsela:'{3, 4, 5, 6, 0, 1, 2}};
  addr_tab[1][1][8][0] = '{baddr:62, offset:'{0, 0, 0, 2047, 2047, 2047, 2047}, offsetm:'{0, 0, 0, 2047, 2047, 2047, 2047}, sela:'{3, 4, 5, 6, 0, 1, 2}, invsela:'{4, 5, 6, 0, 1, 2, 3}};
  addr_tab[1][1][9][0] = '{baddr:65, offset:'{0, 0, 0, 2047, 2047, 2047, 2047}, offsetm:'{0, 0, 0, 2047, 2047, 2047, 2047}, sela:'{3, 4, 5, 6, 0, 1, 2}, invsela:'{4, 5, 6, 0, 1, 2, 3}};
  addr_tab[1][1][10][0] = '{baddr:55, offset:'{0, 2047, 2047, 2047, 2047, 2047, 2047}, offsetm:'{0, 2047, 2047, 2047, 2047, 2047, 2047}, sela:'{1, 2, 3, 4, 5, 6, 0}, invsela:'{6, 0, 1, 2, 3, 4, 5}};
  addr_tab[1][1][11][0] = '{baddr:56, offset:'{0, 2047, 2047, 2047, 2047, 2047, 2047}, offsetm:'{0, 2047, 2047, 2047, 2047, 2047, 2047}, sela:'{1, 2, 3, 4, 5, 6, 0}, invsela:'{6, 0, 1, 2, 3, 4, 5}};
  addr_tab[1][1][12][0] = '{baddr:67, offset:'{0, 0, 0, 0, 0, 2047, 2047}, offsetm:'{0, 0, 0, 0, 0, 2047, 2047}, sela:'{5, 6, 0, 1, 2, 3, 4}, invsela:'{2, 3, 4, 5, 6, 0, 1}};
  addr_tab[1][1][13][0] = '{baddr:68, offset:'{0, 2047, 2047, 2047, 2047, 2047, 2047}, offsetm:'{0, 2047, 2047, 2047, 2047, 2047, 2047}, sela:'{1, 2, 3, 4, 5, 6, 0}, invsela:'{6, 0, 1, 2, 3, 4, 5}};
  addr_tab[1][1][14][0] = '{baddr:55, offset:'{0, 0, 0, 0, 2047, 2047, 2047}, offsetm:'{0, 0, 0, 0, 2047, 2047, 2047}, sela:'{4, 5, 6, 0, 1, 2, 3}, invsela:'{3, 4, 5, 6, 0, 1, 2}};
  addr_tab[1][1][15][0] = '{baddr:60, offset:'{0, 2047, 2047, 2047, 2047, 2047, 2047}, offsetm:'{0, 2047, 2047, 2047, 2047, 2047, 2047}, sela:'{1, 2, 3, 4, 5, 6, 0}, invsela:'{6, 0, 1, 2, 3, 4, 5}};
