localparam int          cLARGE_HS_TAB_1BY4_PACKED_SIZE = 270;
localparam bit [17 : 0] cLARGE_HS_TAB_1BY4_PACKED[cLARGE_HS_TAB_1BY4_PACKED_SIZE] = '{
{1'b0,   8'd0,   9'd4},{1'b1,  8'd27,  9'd69},
{1'b0,  8'd28, 9'd267},{1'b1,  8'd44, 9'd243},
{1'b0,   8'd6,  9'd14},{1'b1,  8'd14,  9'd20},
{1'b0,  8'd13, 9'd332},{1'b1,  8'd20, 9'd325},
{1'b0,   8'd1, 9'd123},{1'b1,  8'd11, 9'd355},
{1'b0,   8'd4, 9'd201},{1'b1,  8'd25, 9'd325},
{1'b0,   8'd5, 9'd103},{1'b1,   8'd5, 9'd189},
{1'b0,  8'd10, 9'd101},{1'b1,  8'd12, 9'd311},
{1'b0,  8'd24, 9'd286},{1'b1,  8'd35, 9'd226},
{1'b0,  8'd17,  9'd47},{1'b1,  8'd41, 9'd219},
{1'b0,   8'd9, 9'd312},{1'b1,  8'd10,  9'd63},
{1'b0,   8'd2,  9'd97},{1'b1,  8'd12,  9'd62},
{1'b0,   8'd8, 9'd223},{1'b1,  8'd15, 9'd164},
{1'b0,  8'd14, 9'd237},{1'b1,  8'd42, 9'd243},
{1'b0,  8'd11, 9'd144},{1'b1,  8'd29,  9'd54},
{1'b0,   8'd0, 9'd137},{1'b1,   8'd2, 9'd224},
{1'b0,   8'd0,  9'd46},{1'b1,   8'd7, 9'd328},
{1'b0,   8'd8, 9'd324},{1'b1,  8'd12,  9'd92},
{1'b0,   8'd9, 9'd206},{1'b1,  8'd40, 9'd126},
{1'b0,   8'd8, 9'd309},{1'b1,  8'd12, 9'd195},
{1'b0,  8'd11, 9'd326},{1'b1,  8'd30,  9'd96},
{1'b0,  8'd14, 9'd203},{1'b1,  8'd23, 9'd179},
{1'b0,   8'd1, 9'd185},{1'b1,  8'd35, 9'd273},
{1'b0,  8'd10, 9'd192},{1'b1,  8'd36,  9'd56},
{1'b0,   8'd6, 9'd333},{1'b1,   8'd8, 9'd214},
{1'b0,   8'd5, 9'd166},{1'b1,  8'd13, 9'd277},
{1'b0,  8'd17, 9'd259},{1'b1,  8'd34, 9'd181},
{1'b0,   8'd3,  9'd66},{1'b1,   8'd4, 9'd213},
{1'b0,   8'd7, 9'd298},{1'b1,  8'd14, 9'd287},
{1'b0,   8'd0, 9'd311},{1'b1,   8'd2, 9'd107},
{1'b0,   8'd6, 9'd312},{1'b1,  8'd30, 9'd125},
{1'b0,   8'd4,  9'd74},{1'b1,   8'd5, 9'd242},
{1'b0,  8'd24, 9'd229},{1'b1,  8'd36, 9'd180},
{1'b0,  8'd11, 9'd180},{1'b1,  8'd25, 9'd263},
{1'b0,   8'd1, 9'd274},{1'b1,   8'd8, 9'd160},
{1'b0,  8'd10, 9'd229},{1'b1,  8'd40,  9'd69},
{1'b0,   8'd4, 9'd299},{1'b1,   8'd6, 9'd171},
{1'b0,   8'd1, 9'd153},{1'b1,   8'd9, 9'd253},
{1'b0,   8'd3, 9'd296},{1'b1,  8'd27, 9'd162},
{1'b0,   8'd9,  9'd33},{1'b1,  8'd19, 9'd106},
{1'b0,   8'd5, 9'd300},{1'b1,  8'd33,  9'd65},
{1'b0,  8'd13, 9'd173},{1'b1,  8'd13, 9'd100},
{1'b0,   8'd0, 9'd176},{1'b1,  8'd16, 9'd143},
{1'b0,  8'd21,  9'd63},{1'b1,  8'd37,   9'd3},
{1'b0,   8'd2,  9'd85},{1'b1,   8'd9,  9'd28},
{1'b0,   8'd5, 9'd136},{1'b1,   8'd8, 9'd155},
{1'b0,   8'd6,  9'd37},{1'b1,  8'd12, 9'd202},
{1'b0,   8'd7, 9'd102},{1'b1,  8'd19, 9'd359},
{1'b0,   8'd6,  9'd76},{1'b1,  8'd11, 9'd126},
{1'b0,  8'd11, 9'd143},{1'b1,  8'd13, 9'd344},
{1'b0,   8'd4, 9'd100},{1'b1,  8'd31, 9'd166},
{1'b0,   8'd7, 9'd278},{1'b1,  8'd13,  9'd23},
{1'b0,   8'd4, 9'd310},{1'b1,   8'd8,  9'd84},
{1'b0,   8'd0, 9'd267},{1'b1,  8'd13, 9'd262},
{1'b0,  8'd11, 9'd112},{1'b1,  8'd23, 9'd151},
{1'b0,   8'd2, 9'd230},{1'b1,  8'd22, 9'd177},
{1'b0,  8'd22, 9'd213},{1'b1,  8'd37, 9'd200},
{1'b0,   8'd6,  9'd65},{1'b1,   8'd9, 9'd281},
{1'b0,   8'd0, 9'd134},{1'b1,  8'd38, 9'd232},
{1'b0,   8'd2, 9'd286},{1'b1,   8'd3,  9'd45},
{1'b0,   8'd0,   9'd8},{1'b1,   8'd7,  9'd88},
{1'b0,  8'd11,  9'd31},{1'b1,  8'd39,  9'd16},
{1'b0,   8'd1, 9'd315},{1'b1,  8'd15,  9'd61},
{1'b0,  8'd14, 9'd317},{1'b1,  8'd41, 9'd128},
{1'b0,   8'd3, 9'd300},{1'b1,  8'd13,  9'd66},
{1'b0,   8'd6, 9'd117},{1'b1,  8'd11, 9'd319},
{1'b0,  8'd13,  9'd43},{1'b1,  8'd33, 9'd350},
{1'b0,   8'd8,  9'd48},{1'b1,  8'd12, 9'd135},
{1'b0,  8'd11,  9'd35},{1'b1,  8'd38,  9'd89},
{1'b0,   8'd9,  9'd42},{1'b1,  8'd35,   9'd6},
{1'b0,   8'd8, 9'd208},{1'b1,  8'd38, 9'd160},
{1'b0,   8'd2, 9'd213},{1'b1,  8'd26,  9'd52},
{1'b0,   8'd4,  9'd59},{1'b1,  8'd34, 9'd111},
{1'b0,   8'd5, 9'd290},{1'b1,   8'd7,  9'd77},
{1'b0,   8'd2, 9'd138},{1'b1,   8'd4,  9'd98},
{1'b0,   8'd9, 9'd201},{1'b1,  8'd10, 9'd290},
{1'b0,  8'd12, 9'd344},{1'b1,  8'd39, 9'd133},
{1'b0,   8'd5,  9'd92},{1'b1,  8'd12, 9'd219},
{1'b0,  8'd14, 9'd285},{1'b1,  8'd26, 9'd111},
{1'b0,  8'd11, 9'd140},{1'b1,  8'd39,   9'd8},
{1'b0,   8'd4, 9'd340},{1'b1,   8'd6, 9'd338},
{1'b0,  8'd11, 9'd218},{1'b1,  8'd17, 9'd248},
{1'b0,  8'd18, 9'd220},{1'b1,  8'd32,  9'd73},
{1'b0,   8'd3, 9'd115},{1'b1,   8'd5, 9'd329},
{1'b0,   8'd1, 9'd121},{1'b1,  8'd31, 9'd175},
{1'b0,   8'd8,   9'd6},{1'b1,  8'd32, 9'd329},
{1'b0,   8'd4, 9'd144},{1'b1,   8'd8, 9'd190},
{1'b0,   8'd7, 9'd243},{1'b1,  8'd24,  9'd60},
{1'b0,   8'd1, 9'd184},{1'b1,   8'd2, 9'd165},
{1'b0,   8'd0, 9'd154},{1'b1,  8'd12, 9'd123},
{1'b0,   8'd8,  9'd49},{1'b1,  8'd12,  9'd69},
{1'b0,   8'd1, 9'd258},{1'b1,  8'd28,  9'd87},
{1'b0,  8'd29, 9'd294},{1'b1,  8'd37,  9'd34},
{1'b0,  8'd18, 9'd218},{1'b1,  8'd42, 9'd341},
{1'b0,   8'd3, 9'd229},{1'b1,  8'd12, 9'd238},
{1'b0,  8'd18, 9'd228},{1'b1,  8'd41, 9'd181},
{1'b0,  8'd12, 9'd262},{1'b1,  8'd15, 9'd179},
{1'b0,  8'd14, 9'd154},{1'b1,  8'd21, 9'd245},
{1'b0,   8'd7, 9'd344},{1'b1,  8'd19,  9'd68},
{1'b0,   8'd2, 9'd103},{1'b1,   8'd9, 9'd264},
{1'b0,   8'd3, 9'd167},{1'b1,  8'd10,  9'd24},
{1'b0,   8'd7,  9'd26},{1'b1,  8'd31,  9'd82},
{1'b0,  8'd13,  9'd53},{1'b1,  8'd44, 9'd152},
{1'b0,   8'd1, 9'd127},{1'b1,  8'd10, 9'd235},
{1'b0,   8'd0, 9'd213},{1'b1,   8'd5, 9'd295},
{1'b0,  8'd27,  9'd40},{1'b1,  8'd40, 9'd286},
{1'b0,  8'd10, 9'd253},{1'b1,  8'd29, 9'd249},
{1'b0,  8'd10,  9'd64},{1'b1,  8'd14, 9'd305},
{1'b0,   8'd0, 9'd348},{1'b1,   8'd6, 9'd335},
{1'b0,   8'd4, 9'd182},{1'b1,  8'd28, 9'd243},
{1'b0,  8'd14, 9'd196},{1'b1,  8'd44, 9'd345},
{1'b0,   8'd6, 9'd143},{1'b1,  8'd10,   9'd8},
{1'b0,  8'd23,  9'd29},{1'b1,  8'd43, 9'd273},
{1'b0,   8'd6, 9'd112},{1'b1,   8'd9,  9'd51},
{1'b0,   8'd3, 9'd164},{1'b1,   8'd3, 9'd124},
{1'b0,   8'd9,  9'd80},{1'b1,  8'd20,  9'd30},
{1'b0,   8'd0, 9'd174},{1'b1,  8'd32, 9'd255},
{1'b0,   8'd1, 9'd155},{1'b1,  8'd13, 9'd115},
{1'b0,   8'd1, 9'd124},{1'b1,  8'd10,  9'd93},
{1'b0,   8'd2,  9'd13},{1'b1,  8'd14,  9'd10},
{1'b0,  8'd21, 9'd254},{1'b1,  8'd43, 9'd135},
{1'b0,  8'd10, 9'd123},{1'b1,  8'd26, 9'd337},
{1'b0,   8'd3, 9'd166},{1'b1,  8'd34, 9'd336},
{1'b0,  8'd16,  9'd73},{1'b1,  8'd43, 9'd150},
{1'b0,   8'd7, 9'd238},{1'b1,  8'd42, 9'd229},
{1'b0,  8'd14, 9'd201},{1'b1,  8'd22, 9'd166},
{1'b0,   8'd4, 9'd242},{1'b1,  8'd20, 9'd281},
{1'b0,  8'd16, 9'd205},{1'b1,  8'd30, 9'd221},
{1'b0,   8'd5, 9'd257},{1'b1,  8'd13, 9'd197},
{1'b0,  8'd14, 9'd347},{1'b1,  8'd25, 9'd158},
{1'b0,   8'd7,  9'd10},{1'b1,  8'd33, 9'd103},
{1'b0,   8'd3,  9'd67},{1'b1,   8'd5,  9'd72},
{1'b0,   8'd3, 9'd176},{1'b1,   8'd9, 9'd162},
{1'b0,   8'd1,  9'd56},{1'b1,   8'd7,  9'd50},
{1'b0,   8'd2, 9'd296},{1'b1,  8'd36,  9'd98}
};
localparam int          cLARGE_HS_TAB_1BY3_PACKED_SIZE = 360;
localparam bit [17 : 0] cLARGE_HS_TAB_1BY3_PACKED[cLARGE_HS_TAB_1BY3_PACKED_SIZE] = '{
{1'b0,   8'd0,  9'd46},{1'b0,   8'd0, 9'd176},{1'b1,  8'd44, 9'd313},
{1'b0,  8'd35, 9'd228},{1'b0,  8'd46, 9'd184},{1'b1,  8'd54, 9'd236},
{1'b0,   8'd6, 9'd143},{1'b0,  8'd16, 9'd243},{1'b1,  8'd27, 9'd284},
{1'b0,   8'd1, 9'd123},{1'b0,  8'd12, 9'd332},{1'b1,  8'd46, 9'd209},
{1'b0,  8'd10, 9'd355},{1'b0,  8'd13,  9'd20},{1'b1,  8'd23, 9'd345},
{1'b0,   8'd4, 9'd201},{1'b0,  8'd17,  9'd86},{1'b1,  8'd18,  9'd16},
{1'b0,   8'd5, 9'd103},{1'b0,   8'd5, 9'd189},{1'b1,  8'd15, 9'd263},
{1'b0,   8'd9, 9'd101},{1'b0,  8'd18, 9'd128},{1'b1,  8'd47,  9'd67},
{1'b0,  8'd21, 9'd145},{1'b0,  8'd22, 9'd133},{1'b1,  8'd34, 9'd330},
{1'b0,   8'd9, 9'd289},{1'b0,  8'd16,  9'd54},{1'b1,  8'd23, 9'd227},
{1'b0,   8'd2,  9'd97},{1'b0,  8'd19, 9'd177},{1'b1,  8'd45, 9'd263},
{1'b0,   8'd8, 9'd312},{1'b0,   8'd9,  9'd63},{1'b1,  8'd16, 9'd108},
{1'b0,  8'd14, 9'd151},{1'b0,  8'd16, 9'd311},{1'b1,  8'd54,  9'd41},
{1'b0,   8'd0, 9'd134},{1'b0,  8'd10, 9'd144},{1'b1,  8'd11,  9'd62},
{1'b0,   8'd0, 9'd137},{1'b0,   8'd2, 9'd224},{1'b1,  8'd22, 9'd323},
{1'b0,   8'd7, 9'd328},{1'b0,  8'd11,  9'd92},{1'b1,  8'd44, 9'd119},
{1'b0,  8'd17,   9'd6},{1'b0,  8'd52,  9'd10},{1'b1,  8'd57,  9'd66},
{1'b0,  8'd13, 9'd237},{1'b0,  8'd34, 9'd176},{1'b1,  8'd35, 9'd245},
{1'b0,   8'd7, 9'd261},{1'b0,   8'd8, 9'd206},{1'b1,  8'd58,  9'd88},
{1'b0,  8'd10, 9'd326},{1'b0,  8'd22, 9'd237},{1'b1,  8'd46, 9'd211},
{1'b0,  8'd10,  9'd97},{1'b0,  8'd14,  9'd63},{1'b1,  8'd32, 9'd332},
{1'b0,   8'd5, 9'd339},{1'b0,  8'd11, 9'd195},{1'b1,  8'd16, 9'd238},
{1'b0,   8'd1, 9'd185},{1'b0,   8'd7, 9'd161},{1'b1,  8'd12, 9'd277},
{1'b0,   8'd3,  9'd66},{1'b0,  8'd17,  9'd73},{1'b1,  8'd29, 9'd148},
{1'b0,   8'd9, 9'd192},{1'b0,  8'd37, 9'd160},{1'b1,  8'd43, 9'd155},
{1'b0,   8'd6,  9'd37},{1'b0,  8'd15, 9'd158},{1'b1,  8'd18, 9'd238},
{1'b0,   8'd0,   9'd4},{1'b0,   8'd5, 9'd166},{1'b1,   8'd8, 9'd254},
{1'b0,   8'd2, 9'd107},{1'b0,   8'd7, 9'd298},{1'b1,  8'd55,  9'd34},
{1'b0,   8'd4, 9'd213},{1'b0,  8'd17,  9'd96},{1'b1,  8'd57, 9'd323},
{1'b0,  8'd13, 9'd187},{1'b0,  8'd20, 9'd235},{1'b1,  8'd41, 9'd214},
{1'b0,   8'd1, 9'd274},{1'b0,   8'd6, 9'd338},{1'b1,  8'd16, 9'd145},
{1'b0,   8'd4, 9'd299},{1'b0,  8'd13, 9'd287},{1'b1,  8'd59, 9'd331},
{1'b0,   8'd5, 9'd242},{1'b0,   8'd6,  9'd14},{1'b1,  8'd19, 9'd315},
{1'b0,  8'd33,   9'd5},{1'b0,  8'd48, 9'd142},{1'b1,  8'd59, 9'd211},
{1'b0,   8'd3, 9'd296},{1'b0,  8'd24, 9'd359},{1'b1,  8'd53, 9'd358},
{1'b0,   8'd5, 9'd300},{1'b0,  8'd15,  9'd57},{1'b1,  8'd15, 9'd139},
{1'b0,  8'd18, 9'd126},{1'b0,  8'd40, 9'd354},{1'b1,  8'd52, 9'd210},
{1'b0,   8'd8, 9'd253},{1'b0,   8'd8,  9'd28},{1'b1,  8'd25, 9'd116},
{1'b0,   8'd0, 9'd154},{1'b0,   8'd6, 9'd335},{1'b1,   8'd9, 9'd229},
{1'b0,  8'd11, 9'd202},{1'b0,  8'd14, 9'd252},{1'b1,  8'd14, 9'd254},
{1'b0,  8'd10, 9'd126},{1'b0,  8'd12, 9'd173},{1'b1,  8'd18,  9'd48},
{1'b0,   8'd2,  9'd85},{1'b0,  8'd16,  9'd14},{1'b1,  8'd53,  9'd72},
{1'b0,   8'd7, 9'd102},{1'b0,  8'd18,  9'd88},{1'b1,  8'd59,  9'd34},
{1'b0,   8'd4, 9'd100},{1'b0,  8'd12,  9'd23},{1'b1,  8'd14, 9'd312},
{1'b0,  8'd18, 9'd181},{1'b0,  8'd30, 9'd332},{1'b1,  8'd48,  9'd82},
{1'b0,   8'd5, 9'd136},{1'b0,  8'd11,  9'd11},{1'b1,  8'd44, 9'd135},
{1'b0,  8'd10, 9'd112},{1'b0,  8'd15, 9'd229},{1'b1,  8'd39,  9'd19},
{1'b0,   8'd0, 9'd174},{1'b0,  8'd17,  9'd56},{1'b1,  8'd50, 9'd123},
{1'b0,  8'd12, 9'd344},{1'b0,  8'd18, 9'd168},{1'b1,  8'd58,  9'd36},
{1'b0,   8'd2, 9'd145},{1'b0,   8'd7, 9'd278},{1'b1,  8'd54, 9'd285},
{1'b0,  8'd12,  9'd66},{1'b0,  8'd16,  9'd87},{1'b1,  8'd18, 9'd101},
{1'b0,   8'd0, 9'd213},{1'b0,  8'd13, 9'd317},{1'b1,  8'd16, 9'd244},
{1'b0,   8'd2, 9'd286},{1'b0,  8'd15,  9'd60},{1'b1,  8'd27,  9'd51},
{1'b0,   8'd0, 9'd267},{1'b0,   8'd4, 9'd310},{1'b1,  8'd19, 9'd212},
{1'b0,  8'd29,  9'd84},{1'b0,  8'd37, 9'd242},{1'b1,  8'd50, 9'd134},
{1'b0,   8'd8, 9'd281},{1'b0,  8'd11, 9'd135},{1'b1,  8'd12,  9'd43},
{1'b0,   8'd1, 9'd315},{1'b0,   8'd3, 9'd300},{1'b1,  8'd43, 9'd327},
{1'b0,   8'd3,  9'd45},{1'b0,   8'd6, 9'd171},{1'b1,  8'd11, 9'd262},
{1'b0,  8'd10,  9'd31},{1'b0,  8'd17, 9'd216},{1'b1,  8'd50, 9'd155},
{1'b0,  8'd20, 9'd207},{1'b0,  8'd25,  9'd41},{1'b1,  8'd36,  9'd24},
{1'b0,   8'd8,  9'd42},{1'b0,  8'd15, 9'd358},{1'b1,  8'd15, 9'd333},
{1'b0,   8'd7,  9'd77},{1'b0,  8'd15, 9'd129},{1'b1,  8'd28, 9'd284},
{1'b0,   8'd2, 9'd213},{1'b0,  8'd17,  9'd58},{1'b1,  8'd53, 9'd206},
{1'b0,   8'd4,  9'd59},{1'b0,   8'd5, 9'd290},{1'b1,  8'd10, 9'd319},
{1'b0,   8'd2, 9'd138},{1'b0,  8'd39, 9'd112},{1'b1,  8'd51, 9'd274},
{1'b0,  8'd10,  9'd35},{1'b0,  8'd23, 9'd228},{1'b1,  8'd29, 9'd122},
{1'b0,   8'd5,  9'd92},{1'b0,  8'd11, 9'd344},{1'b1,  8'd15, 9'd286},
{1'b0,   8'd4,  9'd98},{1'b0,  8'd10, 9'd140},{1'b1,  8'd19, 9'd243},
{1'b0,   8'd8, 9'd201},{1'b0,  8'd11, 9'd123},{1'b1,  8'd56, 9'd120},
{1'b0,  8'd10, 9'd218},{1'b0,  8'd15, 9'd325},{1'b1,  8'd24, 9'd343},
{1'b0,   8'd4, 9'd340},{1'b0,  8'd11, 9'd219},{1'b1,  8'd14, 9'd325},
{1'b0,  8'd17,   9'd3},{1'b0,  8'd18,  9'd69},{1'b1,  8'd32, 9'd242},
{1'b0,   8'd4,  9'd82},{1'b0,  8'd26, 9'd291},{1'b1,  8'd33, 9'd279},
{1'b0,   8'd3, 9'd115},{1'b0,  8'd14,  9'd30},{1'b1,  8'd18, 9'd110},
{1'b0,   8'd1, 9'd121},{1'b0,   8'd6, 9'd333},{1'b1,  8'd11,  9'd69},
{1'b0,   8'd3, 9'd243},{1'b0,  8'd17, 9'd180},{1'b1,  8'd48, 9'd166},
{1'b0,   8'd5, 9'd329},{1'b0,   8'd7, 9'd243},{1'b1,  8'd38, 9'd203},
{1'b0,  8'd37,  9'd44},{1'b0,  8'd38, 9'd238},{1'b1,  8'd56, 9'd184},
{1'b0,   8'd1, 9'd184},{1'b0,   8'd2, 9'd165},{1'b1,  8'd26,  9'd28},
{1'b0,   8'd0, 9'd311},{1'b0,  8'd19, 9'd135},{1'b1,  8'd45, 9'd180},
{1'b0,   8'd4, 9'd144},{1'b0,  8'd14, 9'd120},{1'b1,  8'd27, 9'd239},
{1'b0,   8'd1, 9'd258},{1'b0,  8'd51, 9'd101},{1'b1,  8'd57, 9'd225},
{1'b0,  8'd24,  9'd50},{1'b0,  8'd31,  9'd13},{1'b1,  8'd38,  9'd79},
{1'b0,  8'd11, 9'd238},{1'b0,  8'd13,  9'd44},{1'b1,  8'd13, 9'd154},
{1'b0,  8'd18, 9'd286},{1'b0,  8'd35, 9'd318},{1'b1,  8'd55, 9'd267},
{1'b0,   8'd6, 9'd159},{1'b0,  8'd17, 9'd200},{1'b1,  8'd49, 9'd293},
{1'b0,   8'd9, 9'd192},{1'b0,   8'd9,  9'd24},{1'b1,  8'd19,  9'd61},
{1'b0,  8'd12, 9'd130},{1'b0,  8'd12,  9'd53},{1'b1,  8'd19, 9'd217},
{1'b0,  8'd19, 9'd345},{1'b0,  8'd19,  9'd58},{1'b1,  8'd49, 9'd223},
{1'b0,   8'd2, 9'd103},{1'b0,   8'd3, 9'd167},{1'b1,   8'd9, 9'd235},
{1'b0,  8'd14, 9'd166},{1'b0,  8'd28, 9'd351},{1'b1,  8'd41, 9'd356},
{1'b0,   8'd7,  9'd26},{1'b0,   8'd9, 9'd253},{1'b1,  8'd41, 9'd338},
{1'b0,   8'd0,   9'd8},{1'b0,  8'd14, 9'd168},{1'b1,  8'd36,  9'd84},
{1'b0,   8'd1, 9'd127},{1'b0,  8'd26,  9'd25},{1'b1,  8'd30, 9'd189},
{1'b0,  8'd10, 9'd127},{1'b0,  8'd16, 9'd267},{1'b1,  8'd25, 9'd338},
{1'b0,   8'd5, 9'd295},{1'b0,   8'd8,  9'd51},{1'b1,  8'd31, 9'd121},
{1'b0,   8'd4, 9'd182},{1'b0,   8'd6, 9'd112},{1'b1,  8'd13, 9'd305},
{1'b0,  8'd13,  9'd10},{1'b0,  8'd39, 9'd334},{1'b1,  8'd47,   9'd5},
{1'b0,   8'd6, 9'd117},{1'b0,   8'd9,   9'd8},{1'b1,  8'd42, 9'd267},
{1'b0,   8'd8,  9'd80},{1'b0,  8'd13, 9'd196},{1'b1,  8'd33,  9'd79},
{1'b0,   8'd3, 9'd164},{1'b0,   8'd3, 9'd124},{1'b1,   8'd6, 9'd312},
{1'b0,  8'd28, 9'd341},{1'b0,  8'd32, 9'd308},{1'b1,  8'd45,  9'd56},
{1'b0,   8'd6, 9'd130},{1'b0,  8'd42, 9'd317},{1'b1,  8'd55, 9'd244},
{1'b0,   8'd0, 9'd290},{1'b0,  8'd16, 9'd294},{1'b1,  8'd40, 9'd179},
{1'b0,   8'd1, 9'd155},{1'b0,   8'd8,  9'd95},{1'b1,  8'd56,  9'd21},
{1'b0,   8'd1, 9'd124},{1'b0,   8'd2,  9'd13},{1'b1,   8'd9,  9'd93},
{1'b0,  8'd12, 9'd115},{1'b0,  8'd19, 9'd152},{1'b1,  8'd52, 9'd324},
{1'b0,   8'd9, 9'd123},{1'b0,  8'd12, 9'd103},{1'b1,  8'd43, 9'd348},
{1'b0,  8'd20, 9'd332},{1'b0,  8'd47, 9'd293},{1'b1,  8'd58, 9'd217},
{1'b0,   8'd3, 9'd166},{1'b0,  8'd13, 9'd201},{1'b1,  8'd17, 9'd352},
{1'b0,   8'd7, 9'd238},{1'b0,  8'd15, 9'd107},{1'b1,  8'd49,  9'd69},
{1'b0,  8'd14, 9'd331},{1'b0,  8'd17,  9'd98},{1'b1,  8'd34, 9'd107},
{1'b0,   8'd4, 9'd242},{1'b0,  8'd19, 9'd289},{1'b1,  8'd19, 9'd284},
{1'b0,  8'd16, 9'd332},{1'b0,  8'd21, 9'd324},{1'b1,  8'd31, 9'd129},
{1'b0,  8'd13, 9'd347},{1'b0,  8'd21, 9'd118},{1'b1,  8'd40,  9'd56},
{1'b0,  8'd12, 9'd197},{1'b0,  8'd30, 9'd347},{1'b1,  8'd51,  9'd41},
{1'b0,   8'd1,  9'd96},{1'b0,   8'd5,  9'd72},{1'b1,   8'd7,  9'd10},
{1'b0,   8'd3,  9'd67},{1'b0,   8'd3, 9'd176},{1'b1,  8'd42, 9'd262},
{1'b0,   8'd1,  9'd56},{1'b0,   8'd7,  9'd50},{1'b1,   8'd8, 9'd162},
{1'b0,   8'd2, 9'd296},{1'b0,  8'd14, 9'd245},{1'b1,  8'd36, 9'd303}
};
localparam int          cLARGE_HS_TAB_2BY5_PACKED_SIZE = 432;
localparam bit [17 : 0] cLARGE_HS_TAB_2BY5_PACKED[cLARGE_HS_TAB_2BY5_PACKED_SIZE] = '{
{1'b0,   8'd0,  9'd46},{1'b0,   8'd0, 9'd176},{1'b0,  8'd32, 9'd263},{1'b1,  8'd71, 9'd284},
{1'b0,  8'd17, 9'd243},{1'b0,  8'd19, 9'd128},{1'b0,  8'd23, 9'd173},{1'b1,  8'd45,  9'd66},
{1'b0,   8'd6, 9'd312},{1'b0,  8'd11, 9'd355},{1'b0,  8'd28, 9'd214},{1'b1,  8'd40, 9'd137},
{1'b0,   8'd1, 9'd127},{1'b0,  8'd12, 9'd311},{1'b0,  8'd23, 9'd213},{1'b1,  8'd49, 9'd298},
{1'b0,   8'd5, 9'd189},{1'b0,  8'd13, 9'd332},{1'b0,  8'd16, 9'd263},{1'b1,  8'd71, 9'd137},
{1'b0,   8'd4, 9'd201},{1'b0,   8'd5, 9'd103},{1'b0,  8'd14,  9'd20},{1'b1,  8'd66, 9'd314},
{1'b0,  8'd10, 9'd229},{1'b0,  8'd17,  9'd54},{1'b0,  8'd17, 9'd249},{1'b1,  8'd44, 9'd150},
{1'b0,   8'd9, 9'd312},{1'b0,  8'd24, 9'd160},{1'b0,  8'd32,  9'd61},{1'b1,  8'd61, 9'd317},
{1'b0,   8'd8, 9'd223},{1'b0,  8'd12, 9'd135},{1'b0,  8'd20, 9'd177},{1'b1,  8'd46,  9'd88},
{1'b0,   8'd2,  9'd97},{1'b0,  8'd10,   9'd8},{1'b0,  8'd19, 9'd219},{1'b1,  8'd43, 9'd280},
{1'b0,  8'd11, 9'd144},{1'b0,  8'd18, 9'd226},{1'b0,  8'd21, 9'd230},{1'b1,  8'd67,  9'd99},
{1'b0,  8'd12,  9'd62},{1'b0,  8'd15, 9'd166},{1'b0,  8'd17, 9'd108},{1'b1,  8'd42, 9'd160},
{1'b0,   8'd0, 9'd134},{1'b0,   8'd2, 9'd224},{1'b0,  8'd21,  9'd38},{1'b1,  8'd46, 9'd203},
{1'b0,   8'd0, 9'd137},{1'b0,   8'd7, 9'd328},{1'b0,   8'd8, 9'd309},{1'b1,  8'd60, 9'd205},
{1'b0,  8'd14, 9'd237},{1'b0,  8'd26, 9'd289},{1'b0,  8'd27, 9'd309},{1'b1,  8'd47, 9'd217},
{1'b0,  8'd14, 9'd203},{1'b0,  8'd22, 9'd264},{1'b0,  8'd23, 9'd354},{1'b1,  8'd57, 9'd122},
{1'b0,  8'd15, 9'd245},{1'b0,  8'd17, 9'd238},{1'b0,  8'd21, 9'd186},{1'b1,  8'd59,  9'd97},
{1'b0,   8'd4, 9'd119},{1'b0,   8'd8, 9'd324},{1'b0,  8'd23, 9'd228},{1'b1,  8'd59,  9'd11},
{1'b0,   8'd7, 9'd161},{1'b0,   8'd9, 9'd206},{1'b0,  8'd21, 9'd112},{1'b1,  8'd63, 9'd196},
{1'b0,   8'd6, 9'd335},{1'b0,   8'd8, 9'd214},{1'b0,  8'd11, 9'd326},{1'b1,  8'd68, 9'd122},
{1'b0,   8'd1, 9'd315},{1'b0,   8'd5, 9'd166},{1'b0,  8'd13, 9'd277},{1'b1,  8'd59,  9'd14},
{1'b0,   8'd7, 9'd298},{1'b0,  8'd14, 9'd287},{1'b0,  8'd22,  9'd13},{1'b1,  8'd48, 9'd173},
{1'b0,   8'd2, 9'd107},{1'b0,  8'd12, 9'd195},{1'b0,  8'd16,  9'd52},{1'b1,  8'd56,  9'd70},
{1'b0,   8'd0,   9'd4},{1'b0,   8'd9, 9'd254},{1'b0,  8'd10,  9'd93},{1'b1,  8'd65, 9'd184},
{1'b0,   8'd3,  9'd66},{1'b0,   8'd4,  9'd74},{1'b0,   8'd5, 9'd242},{1'b1,  8'd49, 9'd254},
{1'b0,  8'd16, 9'd158},{1'b0,  8'd19, 9'd126},{1'b0,  8'd24, 9'd176},{1'b1,  8'd56,  9'd98},
{1'b0,   8'd4, 9'd213},{1'b0,   8'd8, 9'd141},{1'b0,  8'd19, 9'd103},{1'b1,  8'd53, 9'd265},
{1'b0,   8'd1, 9'd274},{1'b0,  8'd16,  9'd57},{1'b0,  8'd22, 9'd285},{1'b1,  8'd39, 9'd234},
{1'b0,   8'd6, 9'd333},{1'b0,   8'd8, 9'd160},{1'b0,  8'd34,  9'd75},{1'b1,  8'd50, 9'd279},
{1'b0,   8'd1, 9'd153},{1'b0,   8'd4, 9'd299},{1'b0,  8'd23,  9'd24},{1'b1,  8'd64, 9'd329},
{1'b0,   8'd3, 9'd176},{1'b0,   8'd6, 9'd171},{1'b0,  8'd18, 9'd329},{1'b1,  8'd51, 9'd259},
{1'b0,   8'd6, 9'd143},{1'b0,  8'd11, 9'd180},{1'b0,  8'd27, 9'd354},{1'b1,  8'd53, 9'd182},
{1'b0,   8'd9,  9'd33},{1'b0,  8'd15,  9'd63},{1'b0,  8'd18, 9'd103},{1'b1,  8'd38, 9'd134},
{1'b0,   8'd9, 9'd253},{1'b0,  8'd17, 9'd145},{1'b0,  8'd31, 9'd209},{1'b1,  8'd69, 9'd288},
{1'b0,   8'd0, 9'd154},{1'b0,  8'd10, 9'd192},{1'b0,  8'd15, 9'd312},{1'b1,  8'd57, 9'd248},
{1'b0,   8'd6, 9'd112},{1'b0,  8'd13, 9'd100},{1'b0,  8'd21, 9'd227},{1'b1,  8'd67, 9'd262},
{1'b0,   8'd9,  9'd28},{1'b0,  8'd15, 9'd331},{1'b0,  8'd17,  9'd87},{1'b1,  8'd48, 9'd265},
{1'b0,   8'd2,  9'd85},{1'b0,  8'd11, 9'd126},{1'b0,  8'd33, 9'd271},{1'b1,  8'd65, 9'd107},
{1'b0,   8'd8, 9'd155},{1'b0,  8'd12, 9'd202},{1'b0,  8'd13, 9'd344},{1'b1,  8'd62, 9'd123},
{1'b0,   8'd4, 9'd100},{1'b0,  8'd11, 9'd143},{1'b0,  8'd13, 9'd173},{1'b1,  8'd37,  9'd78},
{1'b0,   8'd7, 9'd102},{1'b0,  8'd16, 9'd139},{1'b0,  8'd22, 9'd121},{1'b1,  8'd50, 9'd293},
{1'b0,   8'd4, 9'd310},{1'b0,   8'd5, 9'd136},{1'b0,  8'd19, 9'd181},{1'b1,  8'd50, 9'd261},
{1'b0,   8'd0, 9'd174},{1'b0,  8'd13, 9'd262},{1'b0,  8'd18, 9'd105},{1'b1,  8'd58, 9'd339},
{1'b0,  8'd11, 9'd112},{1'b0,  8'd18, 9'd255},{1'b0,  8'd25, 9'd294},{1'b1,  8'd68, 9'd202},
{1'b0,   8'd7, 9'd278},{1'b0,  8'd15, 9'd161},{1'b0,  8'd16, 9'd358},{1'b1,  8'd69,  9'd40},
{1'b0,   8'd2, 9'd230},{1'b0,  8'd11,  9'd31},{1'b0,  8'd13,  9'd23},{1'b1,  8'd37, 9'd240},
{1'b0,   8'd0, 9'd213},{1'b0,  8'd23, 9'd318},{1'b0,  8'd32,   9'd9},{1'b1,  8'd58, 9'd147},
{1'b0,   8'd6,  9'd65},{1'b0,  8'd14, 9'd317},{1'b0,  8'd19,  9'd48},{1'b1,  8'd68, 9'd195},
{1'b0,   8'd0, 9'd267},{1'b0,   8'd2, 9'd286},{1'b0,  8'd21, 9'd345},{1'b1,  8'd41,  9'd72},
{1'b0,   8'd3,  9'd67},{1'b0,  8'd11, 9'd319},{1'b0,  8'd20, 9'd315},{1'b1,  8'd37, 9'd123},
{1'b0,   8'd1, 9'd124},{1'b0,   8'd3, 9'd167},{1'b0,  8'd23,  9'd84},{1'b1,  8'd52, 9'd123},
{1'b0,   8'd3, 9'd201},{1'b0,  8'd13,  9'd43},{1'b0,  8'd34, 9'd187},{1'b1,  8'd44,  9'd19},
{1'b0,   8'd9, 9'd281},{1'b0,  8'd12, 9'd344},{1'b0,  8'd27, 9'd230},{1'b1,  8'd69,  9'd44},
{1'b0,  8'd17, 9'd244},{1'b0,  8'd18,  9'd65},{1'b0,  8'd22, 9'd129},{1'b1,  8'd62, 9'd327},
{1'b0,   8'd6,  9'd14},{1'b0,   8'd9,  9'd42},{1'b0,  8'd13,  9'd66},{1'b1,  8'd38, 9'd182},
{1'b0,   8'd8, 9'd208},{1'b0,  8'd18, 9'd350},{1'b0,  8'd19, 9'd168},{1'b1,  8'd57,  9'd96},
{1'b0,   8'd7,  9'd77},{1'b0,   8'd8,  9'd48},{1'b0,  8'd25, 9'd112},{1'b1,  8'd52, 9'd116},
{1'b0,  8'd12, 9'd219},{1'b0,  8'd16, 9'd325},{1'b0,  8'd22, 9'd332},{1'b1,  8'd64, 9'd161},
{1'b0,   8'd2, 9'd138},{1'b0,   8'd2, 9'd213},{1'b0,  8'd10, 9'd290},{1'b1,  8'd47, 9'd312},
{1'b0,   8'd9, 9'd201},{1'b0,  8'd12,  9'd69},{1'b0,  8'd35, 9'd247},{1'b1,  8'd51,  9'd78},
{1'b0,   8'd5, 9'd290},{1'b0,  8'd11,  9'd35},{1'b0,  8'd33, 9'd184},{1'b1,  8'd41,  9'd11},
{1'b0,  8'd11, 9'd140},{1'b0,  8'd14, 9'd285},{1'b0,  8'd20, 9'd212},{1'b1,  8'd46, 9'd359},
{1'b0,   8'd4,  9'd98},{1'b0,   8'd6,  9'd37},{1'b0,  8'd23, 9'd199},{1'b1,  8'd40, 9'd236},
{1'b0,  8'd18, 9'd319},{1'b0,  8'd19, 9'd110},{1'b0,  8'd22, 9'd353},{1'b1,  8'd66, 9'd311},
{1'b0,   8'd4, 9'd340},{1'b0,   8'd5,  9'd92},{1'b0,  8'd19,  9'd69},{1'b1,  8'd45, 9'd181},
{1'b0,   8'd5, 9'd329},{1'b0,  8'd16, 9'd333},{1'b0,  8'd29, 9'd335},{1'b1,  8'd51, 9'd141},
{1'b0,   8'd3, 9'd115},{1'b0,  8'd12, 9'd123},{1'b0,  8'd16, 9'd129},{1'b1,  8'd58, 9'd198},
{1'b0,   8'd1, 9'd184},{1'b0,   8'd8, 9'd190},{1'b0,  8'd30,   9'd1},{1'b1,  8'd36, 9'd275},
{1'b0,   8'd4, 9'd144},{1'b0,  8'd16, 9'd337},{1'b0,  8'd33,  9'd32},{1'b1,  8'd42, 9'd285},
{1'b0,   8'd7, 9'd243},{1'b0,  8'd19, 9'd101},{1'b0,  8'd35, 9'd336},{1'b1,  8'd49, 9'd210},
{1'b0,   8'd1, 9'd123},{1'b0,   8'd8,   9'd6},{1'b0,  8'd19, 9'd329},{1'b1,  8'd42,  9'd49},
{1'b0,   8'd0, 9'd311},{1'b0,  8'd11, 9'd218},{1'b0,  8'd23,  9'd54},{1'b1,  8'd54,  9'd41},
{1'b0,   8'd2, 9'd165},{1'b0,  8'd18, 9'd164},{1'b0,  8'd21, 9'd237},{1'b1,  8'd55, 9'd110},
{1'b0,   8'd1, 9'd155},{1'b0,   8'd8,  9'd49},{1'b0,  8'd20, 9'd243},{1'b1,  8'd43, 9'd250},
{1'b0,  8'd12, 9'd238},{1'b0,  8'd12,  9'd92},{1'b0,  8'd31, 9'd135},{1'b1,  8'd53,  9'd23},
{1'b0,  8'd18,  9'd73},{1'b0,  8'd29,  9'd97},{1'b0,  8'd30,  9'd66},{1'b1,  8'd48, 9'd167},
{1'b0,   8'd3, 9'd229},{1'b0,  8'd15, 9'd252},{1'b0,  8'd24, 9'd252},{1'b1,  8'd38, 9'd340},
{1'b0,  8'd21, 9'd133},{1'b0,  8'd22, 9'd300},{1'b0,  8'd31, 9'd353},{1'b1,  8'd70,  9'd51},
{1'b0,  8'd10,  9'd63},{1'b0,  8'd13,  9'd53},{1'b0,  8'd14, 9'd154},{1'b1,  8'd70,  9'd44},
{1'b0,   8'd3, 9'd166},{1'b0,  8'd12, 9'd262},{1'b0,  8'd18, 9'd349},{1'b1,  8'd71, 9'd156},
{1'b0,   8'd2, 9'd103},{1'b0,   8'd7,  9'd26},{1'b0,   8'd7, 9'd344},{1'b1,  8'd61,  9'd47},
{1'b0,  8'd10,  9'd24},{1'b0,  8'd19, 9'd286},{1'b0,  8'd22,  9'd79},{1'b1,  8'd63,  9'd13},
{1'b0,  8'd20,  9'd61},{1'b0,  8'd20, 9'd217},{1'b0,  8'd23, 9'd303},{1'b1,  8'd39,  9'd67},
{1'b0,   8'd0,   9'd8},{1'b0,   8'd5, 9'd295},{1'b0,  8'd10, 9'd235},{1'b1,  8'd67, 9'd185},
{1'b0,   8'd1,  9'd56},{1'b0,  8'd20, 9'd345},{1'b0,  8'd20,  9'd58},{1'b1,  8'd52, 9'd137},
{1'b0,   8'd6, 9'd130},{1'b0,  8'd10, 9'd253},{1'b0,  8'd18, 9'd200},{1'b1,  8'd65, 9'd306},
{1'b0,  8'd10,  9'd64},{1'b0,  8'd14, 9'd305},{1'b0,  8'd15, 9'd151},{1'b1,  8'd60, 9'd337},
{1'b0,  8'd17, 9'd267},{1'b0,  8'd20, 9'd186},{1'b0,  8'd28, 9'd351},{1'b1,  8'd66,  9'd72},
{1'b0,   8'd4, 9'd182},{1'b0,   8'd9,  9'd51},{1'b0,  8'd26, 9'd112},{1'b1,  8'd36, 9'd125},
{1'b0,   8'd6, 9'd117},{1'b0,  8'd10, 9'd101},{1'b0,  8'd23, 9'd252},{1'b1,  8'd55,  9'd77},
{1'b0,   8'd3, 9'd300},{1'b0,   8'd6, 9'd338},{1'b0,  8'd15, 9'd213},{1'b1,  8'd55, 9'd262},
{1'b0,   8'd3, 9'd124},{1'b0,  8'd14, 9'd196},{1'b0,  8'd30, 9'd327},{1'b1,  8'd36,  9'd69},
{1'b0,   8'd5, 9'd308},{1'b0,   8'd9,  9'd80},{1'b0,  8'd25, 9'd238},{1'b1,  8'd54, 9'd243},
{1'b0,   8'd0, 9'd290},{1'b0,  8'd16, 9'd153},{1'b0,  8'd22, 9'd198},{1'b1,  8'd70,  9'd18},
{1'b0,   8'd1, 9'd258},{1'b0,  8'd13, 9'd115},{1'b0,  8'd20, 9'd152},{1'b1,  8'd45, 9'd296},
{1'b0,   8'd2,  9'd13},{1'b0,  8'd10, 9'd123},{1'b0,  8'd14,  9'd10},{1'b1,  8'd60, 9'd282},
{1'b0,  8'd23, 9'd245},{1'b0,  8'd26, 9'd324},{1'b0,  8'd28, 9'd275},{1'b1,  8'd43, 9'd267},
{1'b0,   8'd3,  9'd45},{1'b0,  8'd20,  9'd81},{1'b0,  8'd21, 9'd194},{1'b1,  8'd56,   9'd8},
{1'b0,   8'd7, 9'd238},{1'b0,  8'd17,  9'd74},{1'b0,  8'd35, 9'd166},{1'b1,  8'd61, 9'd104},
{1'b0,  8'd14, 9'd201},{1'b0,  8'd16, 9'd107},{1'b0,  8'd17, 9'd294},{1'b1,  8'd40, 9'd324},
{1'b0,   8'd4, 9'd242},{1'b0,  8'd15, 9'd177},{1'b0,  8'd29, 9'd317},{1'b1,  8'd39,  9'd41},
{1'b0,  8'd15, 9'd168},{1'b0,  8'd17, 9'd342},{1'b0,  8'd21, 9'd323},{1'b1,  8'd47, 9'd331},
{1'b0,   8'd5, 9'd257},{1'b0,  8'd14, 9'd347},{1'b0,  8'd20, 9'd284},{1'b1,  8'd44, 9'd120},
{1'b0,  8'd13, 9'd197},{1'b0,  8'd21,  9'd27},{1'b0,  8'd21, 9'd228},{1'b1,  8'd54,  9'd57},
{1'b0,   8'd1, 9'd121},{1'b0,   8'd7,  9'd10},{1'b0,  8'd22, 9'd308},{1'b1,  8'd62, 9'd264},
{1'b0,   8'd3, 9'd296},{1'b0,  8'd22, 9'd242},{1'b0,  8'd34, 9'd293},{1'b1,  8'd64, 9'd217},
{1'b0,   8'd1, 9'd185},{1'b0,   8'd5,  9'd72},{1'b0,   8'd9, 9'd162},{1'b1,  8'd63,  9'd82},
{1'b0,   8'd2, 9'd296},{1'b0,   8'd7,  9'd50},{1'b0,  8'd15, 9'd254},{1'b1,  8'd41,   9'd1}
};
localparam int          cLARGE_HS_TAB_1BY2_PACKED_SIZE = 450;
localparam bit [17 : 0] cLARGE_HS_TAB_1BY2_PACKED[cLARGE_HS_TAB_1BY2_PACKED_SIZE] = '{
{1'b0,  8'd26, 9'd300},{1'b0,  8'd27, 9'd259},{1'b0,  8'd30,  9'd67},{1'b0,  8'd36,   9'd0},{1'b1,  8'd74, 9'd181},
{1'b0,  8'd10,  9'd50},{1'b0,  8'd10,  9'd61},{1'b0,  8'd20, 9'd286},{1'b0,  8'd37,   9'd0},{1'b1,  8'd41, 9'd154},
{1'b0,   8'd4,  9'd31},{1'b0,  8'd16,  9'd14},{1'b0,  8'd27, 9'd318},{1'b0,  8'd38,   9'd0},{1'b1,  8'd51, 9'd138},
{1'b0,   8'd2, 9'd262},{1'b0,   8'd6,  9'd69},{1'b0,  8'd16, 9'd267},{1'b0,  8'd39,   9'd0},{1'b1,  8'd68, 9'd352},
{1'b0,   8'd9, 9'd317},{1'b0,  8'd24, 9'd239},{1'b0,  8'd33,  9'd36},{1'b0,  8'd40,   9'd0},{1'b1,  8'd82, 9'd278},
{1'b0,   8'd3, 9'd152},{1'b0,  8'd13, 9'd254},{1'b0,  8'd24, 9'd136},{1'b0,  8'd30, 9'd209},{1'b1,  8'd41,   9'd0},
{1'b0,  8'd14, 9'd286},{1'b0,  8'd21, 9'd103},{1'b0,  8'd32, 9'd236},{1'b0,  8'd42,   9'd0},{1'b1,  8'd76, 9'd338},
{1'b0,   8'd4, 9'd126},{1'b0,  8'd28,  9'd44},{1'b0,  8'd34, 9'd265},{1'b0,  8'd43,   9'd0},{1'b1,  8'd89, 9'd214},
{1'b0,  8'd16, 9'd332},{1'b0,  8'd18,  9'd15},{1'b0,  8'd30, 9'd297},{1'b0,  8'd44,   9'd0},{1'b1,  8'd87,  9'd49},
{1'b0,  8'd21, 9'd341},{1'b0,  8'd24, 9'd341},{1'b0,  8'd45,   9'd0},{1'b0,  8'd58, 9'd296},{1'b1,  8'd79, 9'd353},
{1'b0,   8'd1,  9'd28},{1'b0,   8'd4, 9'd140},{1'b0,   8'd5, 9'd176},{1'b0,  8'd37,   9'd1},{1'b1,  8'd46,   9'd0},
{1'b0,   8'd8, 9'd277},{1'b0,  8'd19, 9'd200},{1'b0,  8'd20, 9'd133},{1'b0,  8'd32, 9'd170},{1'b1,  8'd47,   9'd0},
{1'b0,  8'd15, 9'd333},{1'b0,  8'd26,  9'd79},{1'b0,  8'd33, 9'd181},{1'b0,  8'd48,   9'd0},{1'b1,  8'd78, 9'd197},
{1'b0,   8'd8, 9'd100},{1'b0,  8'd16, 9'd145},{1'b0,  8'd46, 9'd315},{1'b0,  8'd49,   9'd0},{1'b1,  8'd66, 9'd231},
{1'b0,   8'd0,  9'd28},{1'b0,  8'd18, 9'd226},{1'b0,  8'd50,   9'd0},{1'b0,  8'd63, 9'd100},{1'b1,  8'd67, 9'd131},
{1'b0,  8'd13, 9'd166},{1'b0,  8'd23, 9'd335},{1'b0,  8'd30, 9'd184},{1'b0,  8'd51,   9'd0},{1'b1,  8'd63, 9'd299},
{1'b0,   8'd6, 9'd135},{1'b0,  8'd11, 9'd239},{1'b0,  8'd52,   9'd0},{1'b0,  8'd59, 9'd124},{1'b1,  8'd73,  9'd85},
{1'b0,   8'd8, 9'd173},{1'b0,  8'd27,  9'd54},{1'b0,  8'd49, 9'd121},{1'b0,  8'd53,   9'd0},{1'b1,  8'd56, 9'd302},
{1'b0,  8'd14, 9'd110},{1'b0,  8'd23,  9'd51},{1'b0,  8'd25, 9'd273},{1'b0,  8'd54,   9'd0},{1'b1,  8'd81, 9'd161},
{1'b0,   8'd2, 9'd192},{1'b0,  8'd15, 9'd139},{1'b0,  8'd28, 9'd160},{1'b0,  8'd38, 9'd114},{1'b1,  8'd55,   9'd0},
{1'b0,  8'd11,  9'd50},{1'b0,  8'd19,  9'd34},{1'b0,  8'd31, 9'd293},{1'b0,  8'd56,   9'd0},{1'b1,  8'd74,  9'd94},
{1'b0,   8'd0, 9'd306},{1'b0,   8'd8,  9'd23},{1'b0,  8'd11, 9'd188},{1'b0,  8'd57,   9'd0},{1'b1,  8'd67, 9'd280},
{1'b0,  8'd19,  9'd89},{1'b0,  8'd31, 9'd306},{1'b0,  8'd58,   9'd0},{1'b0,  8'd71, 9'd290},{1'b1,  8'd85,  9'd55},
{1'b0,   8'd3, 9'd207},{1'b0,   8'd9,  9'd44},{1'b0,  8'd19, 9'd170},{1'b0,  8'd45, 9'd184},{1'b1,  8'd59,   9'd0},
{1'b0,   8'd4,  9'd35},{1'b0,  8'd17,  9'd73},{1'b0,  8'd35, 9'd204},{1'b0,  8'd52,  9'd97},{1'b1,  8'd60,   9'd0},
{1'b0,  8'd19,   9'd3},{1'b0,  8'd24, 9'd289},{1'b0,  8'd27, 9'd228},{1'b0,  8'd61,   9'd0},{1'b1,  8'd78,  9'd76},
{1'b0,   8'd2, 9'd289},{1'b0,  8'd29, 9'd117},{1'b0,  8'd52,  9'd85},{1'b0,  8'd62,   9'd0},{1'b1,  8'd83, 9'd243},
{1'b0,   8'd7, 9'd130},{1'b0,  8'd13, 9'd168},{1'b0,  8'd34,  9'd69},{1'b0,  8'd63,   9'd0},{1'b1,  8'd66,  9'd19},
{1'b0,  8'd18, 9'd273},{1'b0,  8'd25, 9'd332},{1'b0,  8'd32,  9'd10},{1'b0,  8'd45, 9'd123},{1'b1,  8'd64,   9'd0},
{1'b0,   8'd5, 9'd238},{1'b0,   8'd6, 9'd238},{1'b0,  8'd14,  9'd74},{1'b0,  8'd35, 9'd141},{1'b1,  8'd65,   9'd0},
{1'b0,  8'd20, 9'd126},{1'b0,  8'd22,  9'd61},{1'b0,  8'd47, 9'd155},{1'b0,  8'd66,   9'd0},{1'b1,  8'd86,  9'd30},
{1'b0,   8'd3, 9'd128},{1'b0,   8'd4, 9'd326},{1'b0,  8'd46, 9'd185},{1'b0,  8'd67,   9'd0},{1'b1,  8'd80, 9'd233},
{1'b0,   8'd6, 9'd202},{1'b0,  8'd17, 9'd329},{1'b0,  8'd25, 9'd189},{1'b0,  8'd64, 9'd213},{1'b1,  8'd68,   9'd0},
{1'b0,  8'd15, 9'd111},{1'b0,  8'd16,  9'd87},{1'b0,  8'd35, 9'd293},{1'b0,  8'd40,  9'd46},{1'b1,  8'd69,   9'd0},
{1'b0,  8'd11,  9'd47},{1'b0,  8'd12, 9'd288},{1'b0,  8'd70,   9'd0},{1'b0,  8'd77, 9'd171},{1'b1,  8'd88, 9'd324},
{1'b0,  8'd14, 9'd229},{1'b0,  8'd22, 9'd152},{1'b0,  8'd28, 9'd173},{1'b0,  8'd36, 9'd277},{1'b1,  8'd71,   9'd0},
{1'b0,   8'd5,  9'd35},{1'b0,  8'd21, 9'd229},{1'b0,  8'd25, 9'd277},{1'b0,  8'd51, 9'd296},{1'b1,  8'd72,   9'd0},
{1'b0,   8'd4, 9'd144},{1'b0,  8'd10, 9'd285},{1'b0,  8'd31,  9'd69},{1'b0,  8'd61, 9'd196},{1'b1,  8'd73,   9'd0},
{1'b0,   8'd7, 9'd103},{1'b0,  8'd10, 9'd164},{1'b0,  8'd37,  9'd43},{1'b0,  8'd50,  9'd42},{1'b1,  8'd74,   9'd0},
{1'b0,  8'd20, 9'd101},{1'b0,  8'd26, 9'd332},{1'b0,  8'd48, 9'd357},{1'b0,  8'd55,  9'd95},{1'b1,  8'd75,   9'd0},
{1'b0,  8'd15, 9'd337},{1'b0,  8'd20,  9'd88},{1'b0,  8'd70, 9'd136},{1'b0,  8'd75, 9'd112},{1'b1,  8'd76,   9'd0},
{1'b0,  8'd17, 9'd349},{1'b0,  8'd31, 9'd275},{1'b0,  8'd57, 9'd167},{1'b0,  8'd58,  9'd67},{1'b1,  8'd77,   9'd0},
{1'b0,  8'd16, 9'd311},{1'b0,  8'd20, 9'd238},{1'b0,  8'd27, 9'd245},{1'b0,  8'd78,   9'd0},{1'b1,  8'd86,  9'd73},
{1'b0,  8'd14,  9'd60},{1'b0,  8'd21,  9'd50},{1'b0,  8'd59, 9'd115},{1'b0,  8'd79,   9'd0},{1'b1,  8'd89, 9'd223},
{1'b0,   8'd8,  9'd60},{1'b0,  8'd19, 9'd148},{1'b0,  8'd25, 9'd107},{1'b0,  8'd39,   9'd8},{1'b1,  8'd80,   9'd0},
{1'b0,   8'd1,  9'd51},{1'b0,   8'd5,  9'd68},{1'b0,  8'd18,  9'd58},{1'b0,  8'd22, 9'd177},{1'b1,  8'd81,   9'd0},
{1'b0,   8'd7,  9'd65},{1'b0,  8'd21, 9'd329},{1'b0,  8'd33,  9'd25},{1'b0,  8'd71,  9'd72},{1'b1,  8'd82,   9'd0},
{1'b0,   8'd0,  9'd95},{1'b0,  8'd26, 9'd165},{1'b0,  8'd50, 9'd239},{1'b0,  8'd65, 9'd340},{1'b1,  8'd83,   9'd0},
{1'b0,   8'd0, 9'd103},{1'b0,  8'd10, 9'd179},{1'b0,  8'd14, 9'd204},{1'b0,  8'd35, 9'd211},{1'b1,  8'd84,   9'd0},
{1'b0,   8'd0, 9'd113},{1'b0,   8'd5, 9'd186},{1'b0,  8'd29,  9'd19},{1'b0,  8'd33, 9'd296},{1'b1,  8'd85,   9'd0},
{1'b0,   8'd1, 9'd312},{1'b0,  8'd11, 9'd248},{1'b0,  8'd12, 9'd116},{1'b0,  8'd60, 9'd148},{1'b1,  8'd86,   9'd0},
{1'b0,   8'd1,  9'd40},{1'b0,   8'd3,  9'd64},{1'b0,  8'd21, 9'd243},{1'b0,  8'd85, 9'd229},{1'b1,  8'd87,   9'd0},
{1'b0,   8'd5, 9'd235},{1'b0,  8'd17, 9'd350},{1'b0,  8'd73, 9'd299},{1'b0,  8'd87, 9'd141},{1'b1,  8'd88,   9'd0},
{1'b0,  8'd10, 9'd246},{1'b0,  8'd23, 9'd145},{1'b0,  8'd40, 9'd137},{1'b0,  8'd68, 9'd197},{1'b1,  8'd89,   9'd0},
{1'b0,   8'd0,   9'd0},{1'b0,   8'd3, 9'd290},{1'b0,   8'd6,  9'd92},{1'b0,   8'd8, 9'd262},{1'b1,  8'd83,  9'd50},
{1'b0,   8'd1,   9'd0},{1'b0,  8'd25, 9'd347},{1'b0,  8'd30,   9'd5},{1'b0,  8'd53, 9'd165},{1'b1,  8'd88,   9'd6},
{1'b0,   8'd2,   9'd0},{1'b0,   8'd6, 9'd344},{1'b0,  8'd28, 9'd176},{1'b0,  8'd30,  9'd32},{1'b1,  8'd42,  9'd11},
{1'b0,   8'd3,   9'd0},{1'b0,   8'd3, 9'd171},{1'b0,  8'd12, 9'd106},{1'b0,  8'd26, 9'd308},{1'b1,  8'd60, 9'd106},
{1'b0,   8'd4,   9'd0},{1'b0,   8'd4, 9'd319},{1'b0,  8'd23, 9'd207},{1'b0,  8'd29,  9'd56},{1'b1,  8'd35, 9'd279},
{1'b0,   8'd5,   9'd0},{1'b0,  8'd17, 9'd105},{1'b0,  8'd29, 9'd112},{1'b0,  8'd44,  9'd89},{1'b1,  8'd54, 9'd174},
{1'b0,   8'd6,   9'd0},{1'b0,  8'd12, 9'd359},{1'b0,  8'd21, 9'd311},{1'b0,  8'd38,   9'd2},{1'b1,  8'd57, 9'd300},
{1'b0,   8'd7,   9'd0},{1'b0,  8'd12, 9'd342},{1'b0,  8'd31, 9'd223},{1'b0,  8'd61,  9'd78},{1'b1,  8'd70, 9'd295},
{1'b0,   8'd8,   9'd0},{1'b0,  8'd12,  9'd68},{1'b0,  8'd12,  9'd30},{1'b0,  8'd35,  9'd98},{1'b1,  8'd65, 9'd201},
{1'b0,   8'd1,  9'd80},{1'b0,   8'd1,  9'd33},{1'b0,   8'd9,   9'd0},{1'b0,  8'd29, 9'd324},{1'b1,  8'd34, 9'd132},
{1'b0,   8'd3, 9'd180},{1'b0,  8'd10,   9'd0},{1'b0,  8'd18,  9'd71},{1'b0,  8'd23, 9'd324},{1'b1,  8'd33, 9'd225},
{1'b0,  8'd11,   9'd0},{1'b0,  8'd13, 9'd213},{1'b0,  8'd17, 9'd103},{1'b0,  8'd47, 9'd274},{1'b1,  8'd72, 9'd290},
{1'b0,   8'd7, 9'd253},{1'b0,  8'd12,   9'd0},{1'b0,  8'd15,  9'd52},{1'b0,  8'd24, 9'd351},{1'b1,  8'd81,  9'd77},
{1'b0,   8'd9, 9'd246},{1'b0,  8'd13,   9'd0},{1'b0,  8'd30, 9'd271},{1'b0,  8'd34, 9'd232},{1'b1,  8'd49,  9'd30},
{1'b0,   8'd6, 9'd195},{1'b0,  8'd14,   9'd0},{1'b0,  8'd31, 9'd247},{1'b0,  8'd32, 9'd206},{1'b1,  8'd43,  9'd58},
{1'b0,  8'd15,   9'd0},{1'b0,  8'd22, 9'd345},{1'b0,  8'd26, 9'd126},{1'b0,  8'd79, 9'd138},{1'b1,  8'd84,  9'd88},
{1'b0,   8'd1, 9'd264},{1'b0,  8'd13, 9'd245},{1'b0,  8'd16,   9'd0},{1'b0,  8'd20,  9'd16},{1'b1,  8'd32, 9'd137},
{1'b0,   8'd2, 9'd274},{1'b0,  8'd17,   9'd0},{1'b0,  8'd17, 9'd164},{1'b0,  8'd24, 9'd284},{1'b1,  8'd28,  9'd62},
{1'b0,   8'd2,   9'd8},{1'b0,  8'd18,   9'd0},{1'b0,  8'd34, 9'd173},{1'b0,  8'd39, 9'd267},{1'b1,  8'd53, 9'd224},
{1'b0,  8'd18, 9'd184},{1'b0,  8'd19,   9'd0},{1'b0,  8'd27, 9'd330},{1'b0,  8'd35,  9'd78},{1'b1,  8'd62, 9'd216},
{1'b0,   8'd9, 9'd187},{1'b0,   8'd9, 9'd305},{1'b0,  8'd20,   9'd0},{1'b0,  8'd22, 9'd284},{1'b1,  8'd75, 9'd130},
{1'b0,  8'd21,   9'd0},{1'b0,  8'd22, 9'd217},{1'b0,  8'd23, 9'd352},{1'b0,  8'd69, 9'd103},{1'b1,  8'd77,  9'd14},
{1'b0,  8'd14, 9'd203},{1'b0,  8'd22,   9'd0},{1'b0,  8'd26, 9'd242},{1'b0,  8'd29, 9'd289},{1'b1,  8'd54, 9'd273},
{1'b0,   8'd7, 9'd125},{1'b0,  8'd23,   9'd0},{1'b0,  8'd24, 9'd256},{1'b0,  8'd28, 9'd252},{1'b1,  8'd36, 9'd161},
{1'b0,  8'd13, 9'd151},{1'b0,  8'd15, 9'd275},{1'b0,  8'd24,   9'd0},{1'b0,  8'd41, 9'd176},{1'b1,  8'd44, 9'd312},
{1'b0,   8'd2, 9'd101},{1'b0,  8'd22, 9'd243},{1'b0,  8'd25,   9'd0},{1'b0,  8'd48, 9'd199},{1'b1,  8'd82,  9'd10},
{1'b0,   8'd2,  9'd63},{1'b0,  8'd13, 9'd331},{1'b0,  8'd26,   9'd0},{1'b0,  8'd64,  9'd98},{1'b1,  8'd80, 9'd356},
{1'b0,  8'd16, 9'd243},{1'b0,  8'd27,   9'd0},{1'b0,  8'd34, 9'd253},{1'b0,  8'd72, 9'd124},{1'b1,  8'd76, 9'd333},
{1'b0,   8'd0, 9'd159},{1'b0,   8'd9, 9'd287},{1'b0,  8'd28,   9'd0},{1'b0,  8'd34, 9'd167},{1'b1,  8'd55, 9'd354},
{1'b0,   8'd7, 9'd157},{1'b0,  8'd27,   9'd2},{1'b0,  8'd29,   9'd0},{1'b0,  8'd33, 9'd217},{1'b1,  8'd62,  9'd15},
{1'b0,  8'd11, 9'd189},{1'b0,  8'd18,   9'd6},{1'b0,  8'd28, 9'd242},{1'b0,  8'd30,   9'd0},{1'b1,  8'd69, 9'd329},
{1'b0,   8'd9, 9'd237},{1'b0,  8'd10, 9'd162},{1'b0,  8'd29, 9'd334},{1'b0,  8'd31,   9'd0},{1'b1,  8'd33,  9'd66},
{1'b0,   8'd8, 9'd332},{1'b0,  8'd23, 9'd118},{1'b0,  8'd31, 9'd336},{1'b0,  8'd32,   9'd0},{1'b1,  8'd32, 9'd324},
{1'b0,  8'd11, 9'd259},{1'b0,  8'd25, 9'd353},{1'b0,  8'd33,   9'd0},{1'b0,  8'd42, 9'd236},{1'b1,  8'd84, 9'd241},
{1'b0,   8'd5, 9'd177},{1'b0,   8'd7,   9'd7},{1'b0,  8'd15, 9'd153},{1'b0,  8'd34,   9'd0},{1'b1,  8'd56, 9'd221},
{1'b0,   8'd0, 9'd298},{1'b0,  8'd19, 9'd216},{1'b0,  8'd32, 9'd358},{1'b0,  8'd35,   9'd0},{1'b1,  8'd43, 9'd161}
};
localparam int          cLARGE_HS_TAB_3BY5_PACKED_SIZE = 645;
localparam bit [17 : 0] cLARGE_HS_TAB_3BY5_PACKED[cLARGE_HS_TAB_3BY5_PACKED_SIZE] = '{
{1'b0,   8'd0, 9'd237},{1'b0,  8'd15, 9'd200},{1'b0,  8'd22, 9'd313},{1'b0,  8'd24, 9'd134},{1'b0,  8'd32, 9'd345},{1'b0,  8'd33, 9'd114},{1'b0,  8'd36,   9'd0},{1'b0,  8'd40, 9'd209},{1'b1, 8'd101, 9'd203},
{1'b0,   8'd0, 9'd155},{1'b0,   8'd7, 9'd138},{1'b0,   8'd9,  9'd26},{1'b0,  8'd11, 9'd262},{1'b0,  8'd24,  9'd67},{1'b0,  8'd33, 9'd134},{1'b0,  8'd37,   9'd0},{1'b0,  8'd44,  9'd74},{1'b1,  8'd97, 9'd346},
{1'b0,   8'd2, 9'd357},{1'b0,   8'd6, 9'd257},{1'b0,   8'd8, 9'd178},{1'b0,  8'd14,  9'd52},{1'b0,  8'd33, 9'd156},{1'b0,  8'd34,  9'd35},{1'b0,  8'd38,   9'd0},{1'b0,  8'd64,  9'd94},{1'b1,  8'd92, 9'd339},
{1'b0,  8'd12, 9'd327},{1'b0,  8'd17, 9'd217},{1'b0,  8'd17, 9'd186},{1'b0,  8'd22, 9'd145},{1'b0,  8'd26, 9'd259},{1'b0,  8'd27, 9'd243},{1'b0,  8'd39,   9'd0},{1'b0,  8'd57, 9'd359},{1'b1, 8'd104, 9'd211},
{1'b0,   8'd7, 9'd353},{1'b0,  8'd11, 9'd125},{1'b0,  8'd14, 9'd139},{1'b0,  8'd18,  9'd50},{1'b0,  8'd18, 9'd121},{1'b0,  8'd25,  9'd34},{1'b0,  8'd40,   9'd0},{1'b0,  8'd55,  9'd23},{1'b1,  8'd96, 9'd358},
{1'b0,  8'd22, 9'd209},{1'b0,  8'd24, 9'd210},{1'b0,  8'd25, 9'd160},{1'b0,  8'd28,  9'd11},{1'b0,  8'd29,  9'd53},{1'b0,  8'd31, 9'd120},{1'b0,  8'd41,   9'd0},{1'b0,  8'd48, 9'd201},{1'b1,  8'd94, 9'd137},
{1'b0,   8'd6,  9'd85},{1'b0,  8'd10, 9'd180},{1'b0,  8'd12, 9'd100},{1'b0,  8'd17, 9'd352},{1'b0,  8'd20, 9'd245},{1'b0,  8'd25, 9'd285},{1'b0,  8'd42,   9'd0},{1'b0,  8'd50, 9'd184},{1'b1,  8'd98, 9'd341},
{1'b0,  8'd10,  9'd62},{1'b0,  8'd18, 9'd228},{1'b0,  8'd25, 9'd184},{1'b0,  8'd27, 9'd298},{1'b0,  8'd30,  9'd86},{1'b0,  8'd31,  9'd44},{1'b0,  8'd43,   9'd0},{1'b0,  8'd45, 9'd259},{1'b1,  8'd97, 9'd287},
{1'b0,   8'd3, 9'd354},{1'b0,   8'd8,  9'd88},{1'b0,   8'd8,  9'd98},{1'b0,  8'd22,  9'd56},{1'b0,  8'd35, 9'd246},{1'b0,  8'd38, 9'd130},{1'b0,  8'd44,   9'd0},{1'b1,  8'd79, 9'd357},
{1'b0,   8'd0,  9'd78},{1'b0,   8'd7, 9'd117},{1'b0,  8'd11, 9'd157},{1'b0,  8'd22,  9'd66},{1'b0,  8'd30, 9'd329},{1'b0,  8'd31, 9'd169},{1'b0,  8'd45,   9'd0},{1'b0,  8'd67,  9'd64},{1'b1,  8'd77, 9'd342},
{1'b0,   8'd1,  9'd58},{1'b0,  8'd13,  9'd61},{1'b0,  8'd17,  9'd81},{1'b0,  8'd23, 9'd187},{1'b0,  8'd24, 9'd234},{1'b0,  8'd30, 9'd131},{1'b0,  8'd46,   9'd0},{1'b0,  8'd51, 9'd267},{1'b1, 8'd103,  9'd13},
{1'b0,   8'd4, 9'd106},{1'b0,   8'd9, 9'd300},{1'b0,  8'd11,  9'd92},{1'b0,  8'd11, 9'd136},{1'b0,  8'd15, 9'd336},{1'b0,  8'd16, 9'd243},{1'b0,  8'd47,   9'd0},{1'b0,  8'd56,  9'd61},{1'b1,  8'd82, 9'd288},
{1'b0,   8'd5,  9'd74},{1'b0,  8'd11, 9'd202},{1'b0,  8'd13, 9'd162},{1'b0,  8'd25, 9'd280},{1'b0,  8'd33, 9'd346},{1'b0,  8'd35, 9'd103},{1'b0,  8'd41, 9'd256},{1'b0,  8'd48,   9'd0},{1'b1,  8'd94, 9'd114},
{1'b0,   8'd3,  9'd95},{1'b0,   8'd3, 9'd221},{1'b0,   8'd7,  9'd51},{1'b0,  8'd15, 9'd319},{1'b0,  8'd31,  9'd40},{1'b0,  8'd34, 9'd163},{1'b0,  8'd36, 9'd259},{1'b0,  8'd49,   9'd0},{1'b1,  8'd81,  9'd14},
{1'b0,   8'd7,  9'd65},{1'b0,  8'd13, 9'd285},{1'b0,  8'd15, 9'd111},{1'b0,  8'd17, 9'd332},{1'b0,  8'd28, 9'd318},{1'b0,  8'd29, 9'd352},{1'b0,  8'd50,   9'd0},{1'b0,  8'd69,  9'd28},{1'b1,  8'd89,  9'd96},
{1'b0,   8'd4, 9'd201},{1'b0,  8'd15, 9'd105},{1'b0,  8'd23, 9'd306},{1'b0,  8'd27, 9'd226},{1'b0,  8'd31, 9'd143},{1'b0,  8'd32, 9'd117},{1'b0,  8'd51,   9'd0},{1'b0,  8'd60, 9'd223},{1'b1,  8'd80, 9'd167},
{1'b0,   8'd9, 9'd321},{1'b0,  8'd13, 9'd246},{1'b0,  8'd15,  9'd71},{1'b0,  8'd19, 9'd256},{1'b0,  8'd27, 9'd262},{1'b0,  8'd29,  9'd70},{1'b0,  8'd41, 9'd342},{1'b0,  8'd52,   9'd0},{1'b1, 8'd102,  9'd51},
{1'b0,   8'd2,  9'd30},{1'b0,   8'd5, 9'd352},{1'b0,  8'd23,   9'd5},{1'b0,  8'd26, 9'd204},{1'b0,  8'd29, 9'd319},{1'b0,  8'd35,  9'd88},{1'b0,  8'd53,   9'd0},{1'b0,  8'd60, 9'd300},{1'b1,  8'd90,  9'd86},
{1'b0,   8'd1, 9'd225},{1'b0,   8'd4, 9'd242},{1'b0,  8'd14, 9'd129},{1'b0,  8'd14,  9'd40},{1'b0,  8'd20,  9'd84},{1'b0,  8'd23, 9'd336},{1'b0,  8'd54,   9'd0},{1'b0,  8'd58, 9'd316},{1'b1,  8'd99, 9'd172},
{1'b0,   8'd2, 9'd188},{1'b0,   8'd5,  9'd78},{1'b0,   8'd7, 9'd356},{1'b0,   8'd9, 9'd104},{1'b0,  8'd27,  9'd41},{1'b0,  8'd31,  9'd51},{1'b0,  8'd55,   9'd0},{1'b0,  8'd59, 9'd196},{1'b1,  8'd91, 9'd193},
{1'b0,   8'd2, 9'd121},{1'b0,  8'd10, 9'd290},{1'b0,  8'd11, 9'd307},{1'b0,  8'd19, 9'd122},{1'b0,  8'd23, 9'd166},{1'b0,  8'd32, 9'd304},{1'b0,  8'd56,   9'd0},{1'b0,  8'd63, 9'd112},{1'b1,  8'd92, 9'd183},
{1'b0,   8'd2, 9'd267},{1'b0,   8'd3, 9'd230},{1'b0,   8'd4, 9'd336},{1'b0,   8'd6,  9'd75},{1'b0,  8'd15, 9'd181},{1'b0,  8'd18, 9'd227},{1'b0,  8'd57,   9'd0},{1'b0,  8'd62,   9'd8},{1'b1,  8'd75,  9'd71},
{1'b0,   8'd3, 9'd302},{1'b0,  8'd17,  9'd58},{1'b0,  8'd21, 9'd230},{1'b0,  8'd26, 9'd211},{1'b0,  8'd26, 9'd141},{1'b0,  8'd29, 9'd264},{1'b0,  8'd49,  9'd10},{1'b0,  8'd58,   9'd0},{1'b1, 8'd102, 9'd236},
{1'b0,   8'd1, 9'd236},{1'b0,   8'd9, 9'd285},{1'b0,  8'd19, 9'd289},{1'b0,  8'd27,  9'd57},{1'b0,  8'd27, 9'd110},{1'b0,  8'd42, 9'd266},{1'b0,  8'd59,   9'd0},{1'b1,  8'd79, 9'd304},
{1'b0,   8'd1, 9'd356},{1'b0,   8'd6, 9'd124},{1'b0,  8'd20,  9'd62},{1'b0,  8'd21, 9'd338},{1'b0,  8'd30, 9'd306},{1'b0,  8'd35,  9'd34},{1'b0,  8'd60,   9'd0},{1'b0,  8'd62, 9'd277},{1'b1,  8'd86,  9'd90},
{1'b0,   8'd1, 9'd278},{1'b0,   8'd1, 9'd240},{1'b0,  8'd11, 9'd176},{1'b0,  8'd17, 9'd207},{1'b0,  8'd25,  9'd49},{1'b0,  8'd32, 9'd284},{1'b0,  8'd51, 9'd184},{1'b0,  8'd61,   9'd0},{1'b1,  8'd76, 9'd315},
{1'b0,   8'd0,  9'd43},{1'b0,  8'd14, 9'd275},{1'b0,  8'd16,  9'd48},{1'b0,  8'd17, 9'd212},{1'b0,  8'd28, 9'd284},{1'b0,  8'd35,  9'd21},{1'b0,  8'd52, 9'd293},{1'b0,  8'd62,   9'd0},{1'b1,  8'd76,  9'd96},
{1'b0,   8'd0,   9'd1},{1'b0,   8'd6, 9'd181},{1'b0,  8'd10, 9'd207},{1'b0,  8'd16, 9'd181},{1'b0,  8'd32,  9'd51},{1'b0,  8'd35,  9'd50},{1'b0,  8'd43, 9'd152},{1'b0,  8'd63,   9'd0},{1'b1,  8'd83, 9'd211},
{1'b0,   8'd2,  9'd76},{1'b0,  8'd10,  9'd64},{1'b0,  8'd10, 9'd171},{1'b0,  8'd18, 9'd133},{1'b0,  8'd30, 9'd314},{1'b0,  8'd32, 9'd253},{1'b0,  8'd47, 9'd101},{1'b0,  8'd64,   9'd0},{1'b1,  8'd72, 9'd347},
{1'b0,   8'd2, 9'd317},{1'b0,   8'd5, 9'd280},{1'b0,  8'd10, 9'd228},{1'b0,  8'd11, 9'd311},{1'b0,  8'd27,  9'd94},{1'b0,  8'd30, 9'd228},{1'b0,  8'd59, 9'd149},{1'b0,  8'd65,   9'd0},{1'b1,  8'd75, 9'd294},
{1'b0,   8'd0, 9'd311},{1'b0,   8'd8, 9'd241},{1'b0,   8'd8,  9'd73},{1'b0,  8'd13, 9'd203},{1'b0,  8'd22, 9'd353},{1'b0,  8'd29, 9'd329},{1'b0,  8'd53, 9'd316},{1'b0,  8'd66,   9'd0},{1'b1,  8'd99,  9'd51},
{1'b0,   8'd1, 9'd348},{1'b0,   8'd4, 9'd154},{1'b0,  8'd10, 9'd128},{1'b0,  8'd26, 9'd279},{1'b0,  8'd32,  9'd75},{1'b0,  8'd33, 9'd150},{1'b0,  8'd52,  9'd84},{1'b0,  8'd67,   9'd0},{1'b1,  8'd85, 9'd199},
{1'b0,   8'd6, 9'd290},{1'b0,   8'd7, 9'd197},{1'b0,  8'd21,  9'd19},{1'b0,  8'd22, 9'd135},{1'b0,  8'd23, 9'd142},{1'b0,  8'd32, 9'd223},{1'b0,  8'd66, 9'd188},{1'b0,  8'd68,   9'd0},{1'b1,  8'd88, 9'd122},
{1'b0,   8'd2, 9'd153},{1'b0,   8'd3, 9'd327},{1'b0,   8'd8, 9'd193},{1'b0,  8'd14, 9'd333},{1'b0,  8'd16, 9'd341},{1'b0,  8'd30, 9'd335},{1'b0,  8'd38, 9'd149},{1'b0,  8'd69,   9'd0},{1'b1,  8'd83, 9'd156},
{1'b0,   8'd0, 9'd161},{1'b0,   8'd3,  9'd72},{1'b0,   8'd6,  9'd94},{1'b0,  8'd19, 9'd184},{1'b0,  8'd23, 9'd238},{1'b0,  8'd23,  9'd82},{1'b0,  8'd43, 9'd263},{1'b0,  8'd70,   9'd0},{1'b1, 8'd100, 9'd115},
{1'b0,   8'd0,   9'd2},{1'b0,   8'd3, 9'd174},{1'b0,   8'd3, 9'd160},{1'b0,  8'd13, 9'd164},{1'b0,  8'd24, 9'd331},{1'b0,  8'd27, 9'd324},{1'b0,  8'd36, 9'd257},{1'b0,  8'd71,   9'd0},{1'b1,  8'd96, 9'd241},
{1'b0,   8'd1,  9'd11},{1'b0,   8'd4,  9'd15},{1'b0,   8'd5,  9'd90},{1'b0,  8'd13,  9'd10},{1'b0,  8'd24,  9'd41},{1'b0,  8'd26, 9'd293},{1'b0,  8'd47, 9'd307},{1'b0,  8'd72,   9'd0},{1'b1, 8'd106,  9'd49},
{1'b0,   8'd1, 9'd161},{1'b0,   8'd5, 9'd208},{1'b0,  8'd16, 9'd103},{1'b0,  8'd17, 9'd335},{1'b0,  8'd19, 9'd239},{1'b0,  8'd24, 9'd101},{1'b0,  8'd65,  9'd59},{1'b0,  8'd73,   9'd0},{1'b1, 8'd103, 9'd275},
{1'b0,   8'd9, 9'd319},{1'b0,  8'd11, 9'd253},{1'b0,  8'd12, 9'd277},{1'b0,  8'd25, 9'd324},{1'b0,  8'd34, 9'd266},{1'b0,  8'd35, 9'd192},{1'b0,  8'd44, 9'd277},{1'b0,  8'd74,   9'd0},{1'b1,  8'd74,  9'd68},
{1'b0,  8'd15, 9'd103},{1'b0,  8'd20, 9'd228},{1'b0,  8'd20, 9'd303},{1'b0,  8'd22, 9'd119},{1'b0,  8'd29, 9'd123},{1'b0,  8'd30,  9'd55},{1'b0,  8'd42, 9'd288},{1'b0,  8'd75,   9'd0},{1'b1,  8'd86,  9'd33},
{1'b0,  8'd11, 9'd107},{1'b0,  8'd15,  9'd15},{1'b0,  8'd20, 9'd213},{1'b0,  8'd20, 9'd354},{1'b0,  8'd25,  9'd21},{1'b0,  8'd26,  9'd98},{1'b0,  8'd58, 9'd302},{1'b0,  8'd76,   9'd0},{1'b1, 8'd104, 9'd168},
{1'b0,   8'd4, 9'd229},{1'b0,   8'd9,  9'd40},{1'b0,  8'd25, 9'd267},{1'b0,  8'd25, 9'd341},{1'b0,  8'd30,  9'd72},{1'b0,  8'd34, 9'd346},{1'b0,  8'd49, 9'd154},{1'b0,  8'd77,   9'd0},{1'b1,  8'd93, 9'd187},
{1'b0,   8'd0,  9'd40},{1'b0,   8'd2, 9'd157},{1'b0,  8'd10,  9'd24},{1'b0,  8'd22, 9'd327},{1'b0,  8'd29, 9'd138},{1'b0,  8'd31, 9'd288},{1'b0,  8'd40, 9'd185},{1'b0,  8'd78,   9'd0},{1'b1,  8'd81, 9'd337},
{1'b0,   8'd4, 9'd196},{1'b0,  8'd12,  9'd16},{1'b0,  8'd18, 9'd112},{1'b0,  8'd24, 9'd181},{1'b0,  8'd34, 9'd156},{1'b0,  8'd34,  9'd32},{1'b0,  8'd69, 9'd272},{1'b0,  8'd79,   9'd0},{1'b1,  8'd88, 9'd200},
{1'b0,   8'd8, 9'd298},{1'b0,   8'd8,  9'd55},{1'b0,  8'd12, 9'd173},{1'b0,  8'd15, 9'd350},{1'b0,  8'd20, 9'd199},{1'b0,  8'd26, 9'd273},{1'b0,  8'd64, 9'd132},{1'b0,  8'd80,   9'd0},{1'b1,  8'd82, 9'd194},
{1'b0,   8'd2,  9'd42},{1'b0,   8'd9,  9'd78},{1'b0,  8'd18, 9'd343},{1'b0,  8'd30, 9'd107},{1'b0,  8'd30, 9'd311},{1'b0,  8'd33, 9'd118},{1'b0,  8'd55, 9'd269},{1'b0,  8'd81,   9'd0},{1'b1, 8'd106,  9'd40},
{1'b0,   8'd8, 9'd344},{1'b0,   8'd8,  9'd30},{1'b0,  8'd24, 9'd182},{1'b0,  8'd24, 9'd332},{1'b0,  8'd33,  9'd89},{1'b0,  8'd34,  9'd99},{1'b0,  8'd65, 9'd243},{1'b0,  8'd77, 9'd104},{1'b1,  8'd82,   9'd0},
{1'b0,   8'd7, 9'd125},{1'b0,  8'd13,  9'd50},{1'b0,  8'd21, 9'd324},{1'b0,  8'd26, 9'd261},{1'b0,  8'd26,  9'd78},{1'b0,  8'd35,  9'd39},{1'b0,  8'd54, 9'd274},{1'b0,  8'd83,   9'd0},{1'b1,  8'd91,  9'd56},
{1'b0,   8'd4, 9'd291},{1'b0,  8'd12, 9'd262},{1'b0,  8'd13, 9'd318},{1'b0,  8'd21, 9'd179},{1'b0,  8'd21, 9'd354},{1'b0,  8'd27, 9'd310},{1'b0,  8'd71, 9'd240},{1'b0,  8'd72, 9'd193},{1'b1,  8'd84,   9'd0},
{1'b0,   8'd3, 9'd308},{1'b0,   8'd9, 9'd274},{1'b0,  8'd13, 9'd179},{1'b0,  8'd20,  9'd24},{1'b0,  8'd23, 9'd247},{1'b0,  8'd28,  9'd56},{1'b0,  8'd56,  9'd50},{1'b0,  8'd73, 9'd312},{1'b1,  8'd85,   9'd0},
{1'b0,   8'd5, 9'd131},{1'b0,   8'd7, 9'd233},{1'b0,  8'd14,  9'd11},{1'b0,  8'd20, 9'd252},{1'b0,  8'd29, 9'd327},{1'b0,  8'd32, 9'd137},{1'b0,  8'd37,  9'd41},{1'b0,  8'd86,   9'd0},{1'b1, 8'd107,  9'd47},
{1'b0,   8'd1, 9'd312},{1'b0,  8'd12, 9'd278},{1'b0,  8'd14,  9'd69},{1'b0,  8'd23,  9'd75},{1'b0,  8'd33, 9'd264},{1'b0,  8'd34, 9'd344},{1'b0,  8'd57, 9'd185},{1'b0,  8'd84, 9'd215},{1'b1,  8'd87,   9'd0},
{1'b0,   8'd7,  9'd76},{1'b0,  8'd14, 9'd122},{1'b0,  8'd21, 9'd117},{1'b0,  8'd21,  9'd56},{1'b0,  8'd23, 9'd223},{1'b0,  8'd33, 9'd145},{1'b0,  8'd39, 9'd108},{1'b0,  8'd87, 9'd346},{1'b1,  8'd88,   9'd0},
{1'b0,   8'd0, 9'd277},{1'b0,   8'd7, 9'd330},{1'b0,   8'd9, 9'd312},{1'b0,   8'd9,  9'd33},{1'b0,  8'd13, 9'd114},{1'b0,  8'd28,  9'd68},{1'b0,  8'd61,  9'd51},{1'b0,  8'd78, 9'd177},{1'b1,  8'd89,   9'd0},
{1'b0,  8'd16, 9'd128},{1'b0,  8'd16, 9'd229},{1'b0,  8'd17,  9'd51},{1'b0,  8'd19, 9'd351},{1'b0,  8'd32,  9'd35},{1'b0,  8'd68, 9'd322},{1'b0,  8'd90,   9'd0},{1'b1, 8'd105, 9'd107},
{1'b0,   8'd1,  9'd89},{1'b0,  8'd12, 9'd291},{1'b0,  8'd18, 9'd230},{1'b0,  8'd27, 9'd111},{1'b0,  8'd29, 9'd183},{1'b0,  8'd31, 9'd164},{1'b0,  8'd63,  9'd79},{1'b0,  8'd91,   9'd0},{1'b1, 8'd101, 9'd278},
{1'b0,  8'd15,  9'd65},{1'b0,  8'd16,  9'd50},{1'b0,  8'd18, 9'd345},{1'b0,  8'd18, 9'd359},{1'b0,  8'd22,   9'd1},{1'b0,  8'd22,  9'd25},{1'b0,  8'd68, 9'd161},{1'b0,  8'd92,   9'd0},{1'b1, 8'd105, 9'd316},
{1'b0,   8'd2, 9'd239},{1'b0,   8'd9, 9'd264},{1'b0,  8'd12,  9'd85},{1'b0,  8'd16, 9'd219},{1'b0,  8'd19,  9'd51},{1'b0,  8'd34, 9'd100},{1'b0,  8'd61,  9'd88},{1'b0,  8'd85, 9'd130},{1'b1,  8'd93,   9'd0},
{1'b0,   8'd0, 9'd142},{1'b0,   8'd5,  9'd14},{1'b0,  8'd25, 9'd244},{1'b0,  8'd28, 9'd100},{1'b0,  8'd31, 9'd110},{1'b0,  8'd34,  9'd40},{1'b0,  8'd67,  9'd24},{1'b0,  8'd94,   9'd0},{1'b1,  8'd95,  9'd21},
{1'b0,   8'd3, 9'd352},{1'b0,   8'd4, 9'd148},{1'b0,   8'd5, 9'd197},{1'b0,  8'd12, 9'd332},{1'b0,  8'd16, 9'd329},{1'b0,  8'd19,  9'd70},{1'b0,  8'd39, 9'd170},{1'b0,  8'd74, 9'd174},{1'b1,  8'd95,   9'd0},
{1'b0,   8'd2, 9'd199},{1'b0,   8'd6, 9'd308},{1'b0,  8'd25, 9'd250},{1'b0,  8'd28,  9'd97},{1'b0,  8'd33, 9'd158},{1'b0,  8'd35, 9'd208},{1'b0,  8'd71, 9'd190},{1'b0,  8'd80,  9'd15},{1'b1,  8'd96,   9'd0},
{1'b0,   8'd3, 9'd273},{1'b0,   8'd5, 9'd231},{1'b0,  8'd14, 9'd337},{1'b0,  8'd18, 9'd282},{1'b0,  8'd20, 9'd173},{1'b0,  8'd21, 9'd309},{1'b0,  8'd50, 9'd191},{1'b0,  8'd97,   9'd0},{1'b1, 8'd100,  9'd18},
{1'b0,   8'd0, 9'd114},{1'b0,  8'd12,  9'd60},{1'b0,  8'd29, 9'd296},{1'b0,  8'd30, 9'd184},{1'b0,  8'd32, 9'd156},{1'b0,  8'd33, 9'd227},{1'b0,  8'd37, 9'd145},{1'b0,  8'd84,  9'd64},{1'b1,  8'd98,   9'd0},
{1'b0,   8'd1, 9'd313},{1'b0,   8'd4,  9'd78},{1'b0,  8'd22, 9'd348},{1'b0,  8'd28, 9'd339},{1'b0,  8'd31, 9'd357},{1'b0,  8'd32, 9'd316},{1'b0,  8'd66, 9'd313},{1'b0,  8'd73,  9'd92},{1'b1,  8'd99,   9'd0},
{1'b0,   8'd6,  9'd95},{1'b0,   8'd8, 9'd229},{1'b0,  8'd10, 9'd152},{1'b0,  8'd23, 9'd293},{1'b0,  8'd34, 9'd225},{1'b0,  8'd35, 9'd321},{1'b0,  8'd45, 9'd156},{1'b0,  8'd78, 9'd338},{1'b1, 8'd100,   9'd0},
{1'b0,   8'd7, 9'd273},{1'b0,  8'd14, 9'd153},{1'b0,  8'd17, 9'd235},{1'b0,  8'd26, 9'd194},{1'b0,  8'd31, 9'd236},{1'b0,  8'd35,  9'd82},{1'b0,  8'd70, 9'd188},{1'b0, 8'd101,   9'd0},{1'b1, 8'd107, 9'd107},
{1'b0,   8'd5,  9'd19},{1'b0,  8'd19, 9'd341},{1'b0,  8'd20, 9'd242},{1'b0,  8'd21,  9'd88},{1'b0,  8'd24, 9'd340},{1'b0,  8'd29, 9'd196},{1'b0,  8'd70, 9'd186},{1'b0,  8'd87, 9'd342},{1'b1, 8'd102,   9'd0},
{1'b0,   8'd6, 9'd217},{1'b0,   8'd6, 9'd299},{1'b0,  8'd10,  9'd37},{1'b0,  8'd28, 9'd147},{1'b0,  8'd33,  9'd79},{1'b0,  8'd34, 9'd175},{1'b0,  8'd46, 9'd286},{1'b0,  8'd89,  9'd17},{1'b1, 8'd103,   9'd0},
{1'b0,   8'd4, 9'd216},{1'b0,   8'd5, 9'd119},{1'b0,   8'd6,   9'd6},{1'b0,  8'd14, 9'd111},{1'b0,  8'd17, 9'd315},{1'b0,  8'd26, 9'd173},{1'b0,  8'd53,  9'd80},{1'b0,  8'd95,  9'd83},{1'b1, 8'd104,   9'd0},
{1'b0,  8'd11, 9'd353},{1'b0,  8'd12, 9'd344},{1'b0,  8'd18, 9'd186},{1'b0,  8'd19, 9'd284},{1'b0,  8'd28, 9'd198},{1'b0,  8'd35,   9'd7},{1'b0,  8'd48, 9'd305},{1'b0,  8'd93,  9'd84},{1'b1, 8'd105,   9'd0},
{1'b0,  8'd13, 9'd154},{1'b0,  8'd16, 9'd311},{1'b0,  8'd19, 9'd136},{1'b0,  8'd24, 9'd274},{1'b0,  8'd28,  9'd14},{1'b0,  8'd28,  9'd59},{1'b0,  8'd46, 9'd208},{1'b0,  8'd90, 9'd288},{1'b1, 8'd106,   9'd0},
{1'b0,  8'd10,  9'd10},{1'b0,  8'd15,  9'd76},{1'b0,  8'd19, 9'd196},{1'b0,  8'd21, 9'd112},{1'b0,  8'd21, 9'd289},{1'b0,  8'd31, 9'd341},{1'b0,  8'd54,  9'd58},{1'b0,  8'd98, 9'd285},{1'b1, 8'd107,   9'd0}
};
localparam int          cLARGE_HS_TAB_2BY3_PACKED_SIZE = 480;
localparam bit [17 : 0] cLARGE_HS_TAB_2BY3_PACKED[cLARGE_HS_TAB_2BY3_PACKED_SIZE] = '{
{1'b0,   8'd0,   9'd0},{1'b0,   8'd0,   9'd4},{1'b0,  8'd11, 9'd236},{1'b0,  8'd12, 9'd230},{1'b0,  8'd39, 9'd284},{1'b0,  8'd60,   9'd0},{1'b0,  8'd79, 9'd232},{1'b1,  8'd79, 9'd165},
{1'b0,   8'd1,   9'd0},{1'b0,   8'd3, 9'd189},{1'b0,   8'd7, 9'd311},{1'b0,  8'd12, 9'd236},{1'b0,  8'd17, 9'd225},{1'b0,  8'd61,   9'd0},{1'b0, 8'd111,  9'd61},{1'b1, 8'd112, 9'd302},
{1'b0,   8'd2,   9'd0},{1'b0,   8'd8, 9'd151},{1'b0,  8'd11,  9'd72},{1'b0,  8'd39, 9'd318},{1'b0,  8'd47, 9'd351},{1'b0,  8'd62,   9'd0},{1'b0,  8'd85,  9'd72},{1'b1, 8'd117, 9'd112},
{1'b0,   8'd1, 9'd308},{1'b0,   8'd3,   9'd0},{1'b0,   8'd3, 9'd103},{1'b0,   8'd6, 9'd229},{1'b0,  8'd16,  9'd19},{1'b0,  8'd63,   9'd0},{1'b0, 8'd106, 9'd267},{1'b1, 8'd114, 9'd300},
{1'b0,   8'd1,  9'd97},{1'b0,   8'd2, 9'd201},{1'b0,   8'd4,   9'd0},{1'b0,  8'd30, 9'd339},{1'b0,  8'd58,  9'd31},{1'b0,  8'd64,   9'd0},{1'b0,  8'd72, 9'd266},{1'b1,  8'd78,  9'd34},
{1'b0,   8'd5,   9'd0},{1'b0,   8'd5, 9'd312},{1'b0,   8'd7,  9'd92},{1'b0,   8'd9, 9'd158},{1'b0,  8'd57, 9'd164},{1'b0,  8'd62,  9'd51},{1'b0,  8'd65,   9'd0},{1'b1,  8'd66, 9'd193},
{1'b0,   8'd0, 9'd137},{1'b0,   8'd6,   9'd0},{1'b0,   8'd6,   9'd8},{1'b0,   8'd8, 9'd213},{1'b0,  8'd35,  9'd96},{1'b0,  8'd66,   9'd0},{1'b0,  8'd69,  9'd20},{1'b1,  8'd83, 9'd162},
{1'b0,   8'd0,  9'd46},{1'b0,   8'd1, 9'd224},{1'b0,   8'd7,   9'd0},{1'b0,   8'd7, 9'd344},{1'b0,  8'd14, 9'd267},{1'b0,  8'd67,   9'd0},{1'b0,  8'd88, 9'd123},{1'b1,  8'd99, 9'd286},
{1'b0,   8'd8,   9'd0},{1'b0,  8'd10,   9'd6},{1'b0,  8'd11, 9'd210},{1'b0,  8'd13,  9'd49},{1'b0,  8'd31, 9'd243},{1'b0,  8'd68,   9'd0},{1'b0, 8'd107,  9'd84},{1'b1, 8'd110, 9'd269},
{1'b0,   8'd4, 9'd328},{1'b0,   8'd5, 9'd206},{1'b0,   8'd7, 9'd176},{1'b0,   8'd9,   9'd0},{1'b0,  8'd42, 9'd104},{1'b0,  8'd69,   9'd0},{1'b0,  8'd94,  9'd26},{1'b1, 8'd103, 9'd307},
{1'b0,   8'd6, 9'd207},{1'b0,   8'd7, 9'd135},{1'b0,  8'd10,   9'd0},{1'b0,  8'd38,  9'd68},{1'b0,  8'd42, 9'd317},{1'b0,  8'd70,   9'd0},{1'b0,  8'd85, 9'd133},{1'b1,  8'd94, 9'd125},
{1'b0,   8'd2, 9'd119},{1'b0,   8'd6,  9'd93},{1'b0,   8'd8,  9'd63},{1'b0,  8'd11,   9'd0},{1'b0,  8'd33, 9'd324},{1'b0,  8'd71,   9'd0},{1'b0,  8'd82, 9'd102},{1'b1,  8'd97,   9'd3},
{1'b0,   8'd3, 9'd166},{1'b0,   8'd9, 9'd337},{1'b0,  8'd12,   9'd0},{1'b0,  8'd44, 9'd196},{1'b0,  8'd56,  9'd40},{1'b0,  8'd63, 9'd304},{1'b0,  8'd72,   9'd0},{1'b1, 8'd103, 9'd141},
{1'b0,   8'd0, 9'd311},{1'b0,   8'd1, 9'd107},{1'b0,  8'd11,  9'd67},{1'b0,  8'd13,   9'd0},{1'b0,  8'd40, 9'd337},{1'b0,  8'd65, 9'd169},{1'b0,  8'd73,   9'd0},{1'b1,  8'd76,   9'd4},
{1'b0,   8'd2, 9'd213},{1'b0,   8'd4, 9'd298},{1'b0,  8'd14,   9'd0},{1'b0,  8'd23, 9'd210},{1'b0,  8'd27, 9'd273},{1'b0,  8'd74,   9'd0},{1'b0,  8'd77,  9'd21},{1'b1,  8'd82,  9'd90},
{1'b0,   8'd2,  9'd74},{1'b0,  8'd10,  9'd15},{1'b0,  8'd15,   9'd0},{1'b0,  8'd25, 9'd293},{1'b0,  8'd56, 9'd288},{1'b0,  8'd71, 9'd156},{1'b0,  8'd75,   9'd0},{1'b1, 8'd107, 9'd293},
{1'b0,   8'd3, 9'd242},{1'b0,  8'd10, 9'd226},{1'b0,  8'd16,   9'd0},{1'b0,  8'd19, 9'd359},{1'b0,  8'd34,   9'd8},{1'b0,  8'd76,   9'd0},{1'b0,  8'd86, 9'd260},{1'b1, 8'd102,  9'd84},
{1'b0,   8'd2, 9'd299},{1'b0,   8'd5,  9'd33},{1'b0,   8'd6, 9'd192},{1'b0,  8'd17,   9'd0},{1'b0,  8'd34,  9'd70},{1'b0,  8'd77,   9'd0},{1'b0,  8'd78, 9'd246},{1'b1, 8'd108,  9'd80},
{1'b0,   8'd5, 9'd253},{1'b0,   8'd9, 9'd275},{1'b0,  8'd18,   9'd0},{1'b0,  8'd29, 9'd111},{1'b0,  8'd38,  9'd97},{1'b0,  8'd66, 9'd151},{1'b0,  8'd78,   9'd0},{1'b1,  8'd88, 9'd345},
{1'b0,   8'd0, 9'd176},{1'b0,   8'd9, 9'd333},{1'b0,  8'd19,   9'd0},{1'b0,  8'd47, 9'd196},{1'b0,  8'd50,  9'd55},{1'b0,  8'd67,  9'd89},{1'b0,  8'd79,   9'd0},{1'b1,  8'd84,  9'd91},
{1'b0,   8'd1,  9'd85},{1'b0,   8'd5,  9'd28},{1'b0,  8'd16, 9'd150},{1'b0,  8'd20,   9'd0},{1'b0,  8'd44, 9'd329},{1'b0,  8'd61, 9'd156},{1'b0,  8'd80,   9'd0},{1'b1,  8'd90,  9'd43},
{1'b0,   8'd7, 9'd202},{1'b0,   8'd7, 9'd307},{1'b0,  8'd21,   9'd0},{1'b0,  8'd28, 9'd116},{1'b0,  8'd36, 9'd175},{1'b0,  8'd81,   9'd0},{1'b0,  8'd81, 9'd165},{1'b1,  8'd87, 9'd259},
{1'b0,   8'd3, 9'd136},{1'b0,   8'd8, 9'd161},{1'b0,  8'd22,   9'd0},{1'b0,  8'd48, 9'd161},{1'b0,  8'd55,  9'd86},{1'b0,  8'd70,  9'd18},{1'b0,  8'd74, 9'd133},{1'b1,  8'd82,   9'd0},
{1'b0,   8'd0, 9'd267},{1'b0,   8'd4, 9'd102},{1'b0,  8'd11, 9'd170},{1'b0,  8'd23,   9'd0},{1'b0,  8'd53,  9'd99},{1'b0,  8'd83,   9'd0},{1'b0, 8'd115,  9'd88},{1'b1, 8'd115,  9'd51},
{1'b0,   8'd2, 9'd100},{1'b0,   8'd8, 9'd254},{1'b0,  8'd11, 9'd358},{1'b0,  8'd24,   9'd0},{1'b0,  8'd45, 9'd327},{1'b0,  8'd68, 9'd150},{1'b0,  8'd84,   9'd0},{1'b1,  8'd89, 9'd313},
{1'b0,   8'd0, 9'd134},{1'b0,   8'd1, 9'd230},{1'b0,   8'd9, 9'd325},{1'b0,  8'd25,   9'd0},{1'b0,  8'd37, 9'd198},{1'b0,  8'd85,   9'd0},{1'b0,  8'd98, 9'd311},{1'b1, 8'd105, 9'd272},
{1'b0,   8'd0,   9'd8},{1'b0,   8'd4,  9'd88},{1'b0,  8'd26,   9'd0},{1'b0,  8'd54, 9'd122},{1'b0,  8'd54, 9'd195},{1'b0,  8'd77, 9'd321},{1'b0,  8'd81, 9'd303},{1'b1,  8'd86,   9'd0},
{1'b0,   8'd1, 9'd286},{1'b0,   8'd4, 9'd278},{1'b0,  8'd27,   9'd0},{1'b0,  8'd30, 9'd216},{1'b0,  8'd58, 9'd111},{1'b0,  8'd72, 9'd100},{1'b0,  8'd87,   9'd0},{1'b1,  8'd96, 9'd152},
{1'b0,   8'd2, 9'd310},{1'b0,  8'd10,  9'd76},{1'b0,  8'd10,  9'd58},{1'b0,  8'd22, 9'd167},{1'b0,  8'd28,   9'd0},{1'b0,  8'd88,   9'd0},{1'b0, 8'd105, 9'd212},{1'b1, 8'd113, 9'd149},
{1'b0,   8'd9, 9'd153},{1'b0,  8'd11, 9'd137},{1'b0,  8'd28, 9'd123},{1'b0,  8'd29,   9'd0},{1'b0,  8'd55,  9'd93},{1'b0,  8'd73, 9'd246},{1'b0,  8'd89,   9'd0},{1'b1,  8'd91, 9'd298},
{1'b0,   8'd5, 9'd281},{1'b0,   8'd9, 9'd111},{1'b0,  8'd18,  9'd36},{1'b0,  8'd30,   9'd0},{1'b0,  8'd35, 9'd121},{1'b0,  8'd86,  9'd92},{1'b0,  8'd90,   9'd0},{1'b1,  8'd97, 9'd277},
{1'b0,   8'd4,  9'd77},{1'b0,   8'd6, 9'd290},{1'b0,   8'd7, 9'd238},{1'b0,  8'd11,  9'd10},{1'b0,  8'd31,   9'd0},{1'b0,  8'd91,   9'd0},{1'b0, 8'd100,  9'd56},{1'b1, 8'd117,  9'd79},
{1'b0,   8'd1, 9'd213},{1'b0,   8'd5,  9'd42},{1'b0,   8'd7, 9'd136},{1'b0,  8'd11, 9'd234},{1'b0,  8'd32,   9'd0},{1'b0,  8'd73, 9'd107},{1'b0,  8'd80,   9'd7},{1'b1,  8'd92,   9'd0},
{1'b0,   8'd1, 9'd138},{1'b0,   8'd9, 9'd122},{1'b0,  8'd10, 9'd184},{1'b0,  8'd26,  9'd98},{1'b0,  8'd33,   9'd0},{1'b0,  8'd93,   9'd0},{1'b0, 8'd104, 9'd201},{1'b1, 8'd113, 9'd196},
{1'b0,   8'd3, 9'd290},{1'b0,   8'd7, 9'd195},{1'b0,  8'd34,   9'd0},{1'b0,  8'd52, 9'd131},{1'b0,  8'd57, 9'd341},{1'b0,  8'd65, 9'd178},{1'b0,  8'd69, 9'd272},{1'b1,  8'd94,   9'd0},
{1'b0,   8'd2,  9'd98},{1'b0,  8'd11, 9'd206},{1'b0,  8'd23,   9'd8},{1'b0,  8'd26, 9'd141},{1'b0,  8'd35,   9'd0},{1'b0,  8'd68, 9'd158},{1'b0,  8'd95,   9'd0},{1'b1, 8'd108, 9'd316},
{1'b0,   8'd3,  9'd92},{1'b0,   8'd5, 9'd201},{1'b0,  8'd19, 9'd203},{1'b0,  8'd36,   9'd0},{1'b0,  8'd51,  9'd72},{1'b0,  8'd71, 9'd346},{1'b0,  8'd91, 9'd108},{1'b1,  8'd96,   9'd0},
{1'b0,   8'd2, 9'd340},{1'b0,   8'd3, 9'd329},{1'b0,   8'd9, 9'd129},{1'b0,  8'd20, 9'd331},{1'b0,  8'd37,   9'd0},{1'b0,  8'd97,   9'd0},{1'b0,  8'd98, 9'd259},{1'b1,  8'd99, 9'd348},
{1'b0,   8'd4, 9'd243},{1'b0,   8'd9, 9'd139},{1'b0,  8'd21, 9'd132},{1'b0,  8'd32, 9'd298},{1'b0,  8'd38,   9'd0},{1'b0,  8'd92,   9'd1},{1'b0,  8'd98,   9'd0},{1'b1, 8'd102, 9'd153},
{1'b0,   8'd0, 9'd154},{1'b0,  8'd11, 9'd332},{1'b0,  8'd29, 9'd265},{1'b0,  8'd37, 9'd339},{1'b0,  8'd39,   9'd0},{1'b0,  8'd93, 9'd342},{1'b0,  8'd99,   9'd0},{1'b1, 8'd111,  9'd50},
{1'b0,   8'd1, 9'd165},{1'b0,   8'd7,  9'd69},{1'b0,  8'd22, 9'd265},{1'b0,  8'd40,   9'd0},{1'b0,  8'd53,  9'd72},{1'b0,  8'd95, 9'd266},{1'b0, 8'd100,   9'd0},{1'b1, 8'd118, 9'd132},
{1'b0,   8'd2, 9'd144},{1'b0,   8'd7, 9'd262},{1'b0,  8'd24, 9'd141},{1'b0,  8'd41,   9'd0},{1'b0,  8'd46,  9'd58},{1'b0,  8'd64, 9'd152},{1'b0,  8'd87, 9'd177},{1'b1, 8'd101,   9'd0},
{1'b0,   8'd5, 9'd264},{1'b0,  8'd10, 9'd336},{1'b0,  8'd15, 9'd184},{1'b0,  8'd42,   9'd0},{1'b0,  8'd48, 9'd217},{1'b0,  8'd64, 9'd260},{1'b0,  8'd75, 9'd245},{1'b1, 8'd102,   9'd0},
{1'b0,   8'd6,  9'd24},{1'b0,   8'd9,  9'd52},{1'b0,  8'd27, 9'd173},{1'b0,  8'd33, 9'd111},{1'b0,  8'd43,   9'd0},{1'b0,  8'd96, 9'd171},{1'b0, 8'd103,   9'd0},{1'b1, 8'd109, 9'd274},
{1'b0,   8'd1, 9'd103},{1'b0,   8'd4, 9'd344},{1'b0,  8'd25, 9'd279},{1'b0,  8'd44,   9'd0},{1'b0,  8'd59, 9'd342},{1'b0,  8'd90, 9'd149},{1'b0,  8'd93,  9'd61},{1'b1, 8'd104,   9'd0},
{1'b0,   8'd6, 9'd235},{1'b0,  8'd10, 9'd181},{1'b0,  8'd36, 9'd148},{1'b0,  8'd41, 9'd322},{1'b0,  8'd45,   9'd0},{1'b0,  8'd76,  9'd50},{1'b0,  8'd84, 9'd200},{1'b1, 8'd105,   9'd0},
{1'b0,   8'd0, 9'd213},{1'b0,   8'd8, 9'd320},{1'b0,  8'd15, 9'd341},{1'b0,  8'd41, 9'd325},{1'b0,  8'd46,   9'd0},{1'b0,  8'd60, 9'd303},{1'b0,  8'd61, 9'd137},{1'b1, 8'd106,   9'd0},
{1'b0,   8'd6, 9'd253},{1'b0,   8'd6,  9'd64},{1'b0,  8'd13, 9'd160},{1'b0,  8'd47,   9'd0},{1'b0,  8'd50, 9'd184},{1'b0,  8'd60, 9'd286},{1'b0, 8'd107,   9'd0},{1'b1, 8'd114, 9'd223},
{1'b0,   8'd0, 9'd348},{1'b0,   8'd4,  9'd26},{1'b0,  8'd18,  9'd25},{1'b0,  8'd45, 9'd123},{1'b0,  8'd48,   9'd0},{1'b0,  8'd92, 9'd185},{1'b0, 8'd108,   9'd0},{1'b1, 8'd116, 9'd277},
{1'b0,   8'd3, 9'd295},{1'b0,   8'd5,  9'd51},{1'b0,  8'd10, 9'd111},{1'b0,  8'd21,  9'd69},{1'b0,  8'd49,   9'd0},{1'b0,  8'd75, 9'd234},{1'b0, 8'd109,   9'd0},{1'b1, 8'd119,  9'd59},
{1'b0,   8'd2, 9'd182},{1'b0,   8'd8, 9'd166},{1'b0,  8'd24, 9'd140},{1'b0,  8'd31,  9'd41},{1'b0,  8'd50,   9'd0},{1'b0, 8'd110,   9'd0},{1'b0, 8'd112, 9'd316},{1'b1, 8'd119, 9'd243},
{1'b0,   8'd0, 9'd174},{1'b0,   8'd5,  9'd80},{1'b0,   8'd6, 9'd101},{1'b0,  8'd10, 9'd352},{1'b0,  8'd51,   9'd0},{1'b0,  8'd74, 9'd309},{1'b0, 8'd111,   9'd0},{1'b1, 8'd116,   9'd8},
{1'b0,   8'd3, 9'd308},{1'b0,   8'd8, 9'd168},{1'b0,  8'd40, 9'd205},{1'b0,  8'd51, 9'd314},{1'b0,  8'd52,   9'd0},{1'b0,  8'd95, 9'd194},{1'b0, 8'd101, 9'd334},{1'b1, 8'd112,   9'd0},
{1'b0,   8'd6, 9'd123},{1'b0,  8'd10, 9'd273},{1'b0,  8'd14, 9'd244},{1'b0,  8'd43, 9'd319},{1'b0,  8'd53,   9'd0},{1'b0,  8'd62, 9'd117},{1'b0, 8'd104, 9'd345},{1'b1, 8'd113,   9'd0},
{1'b0,   8'd8,  9'd90},{1'b0,  8'd11, 9'd324},{1'b0,  8'd17,  9'd66},{1'b0,  8'd49, 9'd148},{1'b0,  8'd54,   9'd0},{1'b0,  8'd70, 9'd249},{1'b0,  8'd80, 9'd122},{1'b1, 8'd114,   9'd0},
{1'b0,   8'd4, 9'd238},{1'b0,   8'd8, 9'd177},{1'b0,  8'd20,  9'd34},{1'b0,  8'd32, 9'd110},{1'b0,  8'd55,   9'd0},{1'b0, 8'd106, 9'd184},{1'b0, 8'd115,   9'd0},{1'b1, 8'd118,  9'd94},
{1'b0,   8'd2, 9'd242},{1'b0,   8'd9,  9'd11},{1'b0,  8'd46, 9'd267},{1'b0,  8'd56,   9'd0},{1'b0,  8'd59,  9'd86},{1'b0, 8'd100,  9'd70},{1'b0, 8'd109,  9'd58},{1'b1, 8'd116,   9'd0},
{1'b0,   8'd3, 9'd257},{1'b0,  8'd10,  9'd71},{1'b0,  8'd43, 9'd183},{1'b0,  8'd49,  9'd86},{1'b0,  8'd57,   9'd0},{1'b0,  8'd63, 9'd223},{1'b0,  8'd83, 9'd167},{1'b1, 8'd117,   9'd0},
{1'b0,   8'd4,  9'd50},{1'b0,   8'd5, 9'd162},{1'b0,   8'd8, 9'd331},{1'b0,  8'd52,  9'd64},{1'b0,  8'd58,   9'd0},{1'b0,  8'd67, 9'd156},{1'b0,  8'd89,  9'd41},{1'b1, 8'd118,   9'd0},
{1'b0,   8'd1, 9'd296},{1'b0,   8'd3,  9'd72},{1'b0,   8'd4,  9'd10},{1'b0,   8'd8, 9'd245},{1'b0,  8'd59,   9'd0},{1'b0, 8'd101, 9'd286},{1'b0, 8'd110,  9'd23},{1'b1, 8'd119,   9'd0}
};
localparam int          cLARGE_HS_TAB_3BY4_PACKED_SIZE = 539;
localparam bit [17 : 0] cLARGE_HS_TAB_3BY4_PACKED[cLARGE_HS_TAB_3BY4_PACKED_SIZE] = '{
{1'b0,   8'd0,   9'd0},{1'b0,   8'd2, 9'd308},{1'b0,   8'd3, 9'd155},{1'b0,   8'd6, 9'd215},{1'b0,  8'd10, 9'd196},{1'b0,  8'd31,  9'd97},{1'b0,  8'd45,   9'd0},{1'b0,  8'd59, 9'd187},{1'b0,  8'd69,  9'd59},{1'b0,  8'd90,   9'd0},{1'b0,  8'd94, 9'd173},{1'b1, 8'd126, 9'd282},
{1'b0,   8'd1,   9'd0},{1'b0,   8'd3,  9'd81},{1'b0,   8'd7,   9'd9},{1'b0,   8'd9,  9'd46},{1'b0,  8'd39, 9'd318},{1'b0,  8'd40, 9'd181},{1'b0,  8'd46,   9'd0},{1'b0,  8'd62, 9'd268},{1'b0,  8'd82, 9'd209},{1'b0,  8'd91,   9'd0},{1'b0, 8'd113, 9'd331},{1'b1, 8'd129, 9'd180},
{1'b0,   8'd1, 9'd150},{1'b0,   8'd2,   9'd0},{1'b0,   8'd2, 9'd271},{1'b0,   8'd7, 9'd338},{1'b0,  8'd30,  9'd70},{1'b0,  8'd40, 9'd347},{1'b0,  8'd47,   9'd0},{1'b0,  8'd51, 9'd176},{1'b0,  8'd85, 9'd327},{1'b0,  8'd90, 9'd157},{1'b0,  8'd92,   9'd0},{1'b1, 8'd114, 9'd332},
{1'b0,   8'd3,   9'd0},{1'b0,   8'd5, 9'd140},{1'b0,   8'd7,  9'd88},{1'b0,   8'd8,  9'd12},{1'b0,   8'd8, 9'd309},{1'b0,  8'd17, 9'd291},{1'b0,  8'd48,   9'd0},{1'b0,  8'd48, 9'd262},{1'b0,  8'd50, 9'd155},{1'b0,  8'd93,   9'd0},{1'b0, 8'd123, 9'd165},{1'b1, 8'd134,  9'd64},
{1'b0,   8'd2, 9'd321},{1'b0,   8'd4,   9'd0},{1'b0,  8'd10, 9'd157},{1'b0,  8'd11, 9'd347},{1'b0,  8'd29, 9'd191},{1'b0,  8'd36,  9'd41},{1'b0,  8'd45,  9'd28},{1'b0,  8'd46, 9'd280},{1'b0,  8'd49,   9'd0},{1'b0,  8'd94,   9'd0},{1'b0, 8'd100,  9'd20},{1'b1, 8'd107, 9'd189},
{1'b0,   8'd5,   9'd0},{1'b0,   8'd5, 9'd278},{1'b0,   8'd9, 9'd161},{1'b0,  8'd30,  9'd77},{1'b0,  8'd32, 9'd305},{1'b0,  8'd50,   9'd0},{1'b0,  8'd73, 9'd356},{1'b0,  8'd77, 9'd269},{1'b0,  8'd94,  9'd31},{1'b0,  8'd95,   9'd0},{1'b1, 8'd131, 9'd336},
{1'b0,   8'd5, 9'd315},{1'b0,   8'd6,   9'd0},{1'b0,   8'd8, 9'd204},{1'b0,   8'd9,  9'd12},{1'b0,  8'd12, 9'd194},{1'b0,  8'd16, 9'd298},{1'b0,  8'd48,  9'd70},{1'b0,  8'd51,   9'd0},{1'b0,  8'd89, 9'd138},{1'b0,  8'd96,   9'd0},{1'b0,  8'd98, 9'd107},{1'b1, 8'd106,  9'd61},
{1'b0,   8'd7,   9'd0},{1'b0,   8'd9, 9'd281},{1'b0,  8'd13, 9'd150},{1'b0,  8'd14, 9'd181},{1'b0,  8'd19, 9'd160},{1'b0,  8'd33, 9'd315},{1'b0,  8'd47,  9'd60},{1'b0,  8'd52,   9'd0},{1'b0,  8'd66,  9'd87},{1'b0,  8'd97,   9'd0},{1'b0, 8'd108, 9'd198},{1'b1, 8'd123, 9'd299},
{1'b0,   8'd4,  9'd36},{1'b0,   8'd8,   9'd0},{1'b0,   8'd8,  9'd79},{1'b0,  8'd10, 9'd224},{1'b0,  8'd12, 9'd328},{1'b0,  8'd21,  9'd98},{1'b0,  8'd53,   9'd0},{1'b0,  8'd55,  9'd39},{1'b0,  8'd89, 9'd171},{1'b0,  8'd96, 9'd171},{1'b0,  8'd98,   9'd0},{1'b1, 8'd116, 9'd146},
{1'b0,   8'd1, 9'd307},{1'b0,   8'd2, 9'd142},{1'b0,   8'd4, 9'd240},{1'b0,   8'd6,  9'd90},{1'b0,   8'd9,   9'd0},{1'b0,  8'd29, 9'd285},{1'b0,  8'd54,   9'd0},{1'b0,  8'd57,  9'd12},{1'b0,  8'd87,  9'd26},{1'b0,  8'd99,   9'd0},{1'b0, 8'd108, 9'd271},{1'b1, 8'd111,  9'd89},
{1'b0,   8'd1, 9'd340},{1'b0,   8'd4, 9'd108},{1'b0,   8'd9, 9'd147},{1'b0,  8'd10,   9'd0},{1'b0,  8'd12,  9'd81},{1'b0,  8'd13,  9'd11},{1'b0,  8'd55,   9'd0},{1'b0,  8'd63, 9'd179},{1'b0,  8'd78, 9'd344},{1'b0,  8'd99, 9'd265},{1'b0, 8'd100,   9'd0},{1'b1, 8'd100,  9'd40},
{1'b0,   8'd0,  9'd18},{1'b0,   8'd5, 9'd120},{1'b0,   8'd8, 9'd128},{1'b0,  8'd11,   9'd0},{1'b0,  8'd15, 9'd266},{1'b0,  8'd23, 9'd168},{1'b0,  8'd56,   9'd0},{1'b0,  8'd56,  9'd38},{1'b0,  8'd57, 9'd276},{1'b0,  8'd97,  9'd57},{1'b0, 8'd101,   9'd0},{1'b1, 8'd122, 9'd272},
{1'b0,   8'd0,  9'd72},{1'b0,   8'd2, 9'd177},{1'b0,  8'd12,   9'd0},{1'b0,  8'd12, 9'd109},{1'b0,  8'd13,  9'd58},{1'b0,  8'd31, 9'd309},{1'b0,  8'd52, 9'd335},{1'b0,  8'd57,   9'd0},{1'b0,  8'd76, 9'd213},{1'b0,  8'd90,  9'd77},{1'b0, 8'd102,   9'd0},{1'b1, 8'd104, 9'd174},
{1'b0,   8'd4, 9'd206},{1'b0,  8'd10, 9'd205},{1'b0,  8'd11,  9'd42},{1'b0,  8'd13,   9'd0},{1'b0,  8'd13, 9'd198},{1'b0,  8'd41, 9'd249},{1'b0,  8'd53, 9'd112},{1'b0,  8'd58,   9'd0},{1'b0,  8'd68,  9'd39},{1'b0, 8'd103,   9'd0},{1'b0, 8'd107, 9'd103},{1'b1, 8'd110, 9'd280},
{1'b0,   8'd3, 9'd262},{1'b0,   8'd4, 9'd215},{1'b0,  8'd12, 9'd354},{1'b0,  8'd13, 9'd294},{1'b0,  8'd14,   9'd0},{1'b0,  8'd22,  9'd59},{1'b0,  8'd51, 9'd357},{1'b0,  8'd59,   9'd0},{1'b0,  8'd62,  9'd31},{1'b0, 8'd104,   9'd0},{1'b0, 8'd105, 9'd135},{1'b1, 8'd116, 9'd190},
{1'b0,   8'd4,  9'd27},{1'b0,   8'd7, 9'd267},{1'b0,  8'd10, 9'd146},{1'b0,  8'd15,   9'd0},{1'b0,  8'd18, 9'd321},{1'b0,  8'd26, 9'd136},{1'b0,  8'd60,   9'd0},{1'b0,  8'd68, 9'd130},{1'b0,  8'd86, 9'd341},{1'b0, 8'd102,  9'd79},{1'b0, 8'd105,   9'd0},{1'b1, 8'd125,  9'd56},
{1'b0,   8'd3, 9'd162},{1'b0,   8'd6, 9'd196},{1'b0,   8'd6, 9'd103},{1'b0,   8'd9, 9'd217},{1'b0,  8'd16,   9'd0},{1'b0,  8'd35, 9'd117},{1'b0,  8'd61,   9'd0},{1'b0,  8'd84, 9'd189},{1'b0,  8'd85, 9'd188},{1'b0,  8'd91,  9'd87},{1'b0, 8'd106,   9'd0},{1'b1, 8'd114, 9'd158},
{1'b0,   8'd2, 9'd336},{1'b0,   8'd3, 9'd295},{1'b0,   8'd3, 9'd318},{1'b0,  8'd17,   9'd0},{1'b0,  8'd28, 9'd192},{1'b0,  8'd39, 9'd170},{1'b0,  8'd62,   9'd0},{1'b0,  8'd69, 9'd332},{1'b0,  8'd88,  9'd52},{1'b0, 8'd102, 9'd251},{1'b0, 8'd107,   9'd0},{1'b1, 8'd129, 9'd226},
{1'b0,   8'd6, 9'd230},{1'b0,   8'd6, 9'd228},{1'b0,   8'd7, 9'd203},{1'b0,  8'd11, 9'd240},{1'b0,  8'd14, 9'd321},{1'b0,  8'd18,   9'd0},{1'b0,  8'd50, 9'd312},{1'b0,  8'd60, 9'd217},{1'b0,  8'd63,   9'd0},{1'b0, 8'd108,   9'd0},{1'b0, 8'd119, 9'd308},{1'b1, 8'd121, 9'd255},
{1'b0,   8'd1, 9'd252},{1'b0,   8'd4, 9'd324},{1'b0,  8'd12,  9'd47},{1'b0,  8'd13, 9'd346},{1'b0,  8'd19,   9'd0},{1'b0,  8'd35, 9'd334},{1'b0,  8'd64,   9'd0},{1'b0,  8'd77, 9'd342},{1'b0,  8'd87, 9'd176},{1'b0,  8'd96,  9'd55},{1'b0, 8'd109,   9'd0},{1'b1, 8'd127, 9'd207},
{1'b0,   8'd5, 9'd309},{1'b0,   8'd8,  9'd19},{1'b0,  8'd10, 9'd246},{1'b0,  8'd20,   9'd0},{1'b0,  8'd27, 9'd166},{1'b0,  8'd38, 9'd135},{1'b0,  8'd46, 9'd221},{1'b0,  8'd65,   9'd0},{1'b0,  8'd74, 9'd103},{1'b0, 8'd110,   9'd0},{1'b0, 8'd113,  9'd38},{1'b1, 8'd132, 9'd321},
{1'b0,   8'd1,  9'd44},{1'b0,   8'd2, 9'd140},{1'b0,   8'd4, 9'd169},{1'b0,  8'd11, 9'd245},{1'b0,  8'd16, 9'd153},{1'b0,  8'd21,   9'd0},{1'b0,  8'd56, 9'd180},{1'b0,  8'd66,   9'd0},{1'b0,  8'd82, 9'd106},{1'b0, 8'd103, 9'd331},{1'b0, 8'd110,  9'd98},{1'b1, 8'd111,   9'd0},
{1'b0,   8'd0,  9'd60},{1'b0,   8'd2, 9'd302},{1'b0,   8'd4, 9'd253},{1'b0,   8'd8, 9'd133},{1'b0,   8'd9, 9'd162},{1'b0,  8'd22,   9'd0},{1'b0,  8'd67,   9'd0},{1'b0,  8'd81, 9'd183},{1'b0,  8'd84,  9'd62},{1'b0,  8'd98, 9'd348},{1'b0, 8'd112,   9'd0},{1'b1, 8'd120, 9'd263},
{1'b0,   8'd0, 9'd116},{1'b0,   8'd5, 9'd163},{1'b0,   8'd6, 9'd174},{1'b0,  8'd23,   9'd0},{1'b0,  8'd23, 9'd200},{1'b0,  8'd36,  9'd24},{1'b0,  8'd55, 9'd343},{1'b0,  8'd64, 9'd187},{1'b0,  8'd68,   9'd0},{1'b0, 8'd106,  9'd87},{1'b0, 8'd109, 9'd276},{1'b1, 8'd113,   9'd0},
{1'b0,   8'd0, 9'd297},{1'b0,   8'd9,  9'd75},{1'b0,  8'd11, 9'd328},{1'b0,  8'd24,   9'd0},{1'b0,  8'd27, 9'd323},{1'b0,  8'd38, 9'd214},{1'b0,  8'd69,   9'd0},{1'b0,  8'd78, 9'd194},{1'b0,  8'd80, 9'd345},{1'b0, 8'd114,   9'd0},{1'b0, 8'd124, 9'd291},{1'b1, 8'd133, 9'd247},
{1'b0,   8'd8, 9'd138},{1'b0,   8'd9, 9'd106},{1'b0,  8'd11, 9'd256},{1'b0,  8'd22, 9'd310},{1'b0,  8'd25,   9'd0},{1'b0,  8'd42, 9'd303},{1'b0,  8'd70,   9'd0},{1'b0,  8'd79, 9'd340},{1'b0,  8'd81,  9'd66},{1'b0,  8'd92, 9'd170},{1'b0, 8'd115,   9'd0},{1'b1, 8'd118, 9'd284},
{1'b0,   8'd0, 9'd175},{1'b0,   8'd7, 9'd271},{1'b0,  8'd14,  9'd67},{1'b0,  8'd14, 9'd145},{1'b0,  8'd25, 9'd161},{1'b0,  8'd26,   9'd0},{1'b0,  8'd58, 9'd157},{1'b0,  8'd67,  9'd85},{1'b0,  8'd71,   9'd0},{1'b0, 8'd116,   9'd0},{1'b0, 8'd120, 9'd248},{1'b1, 8'd128, 9'd341},
{1'b0,   8'd6, 9'd177},{1'b0,   8'd8, 9'd315},{1'b0,   8'd9, 9'd109},{1'b0,  8'd20,  9'd73},{1'b0,  8'd27,   9'd0},{1'b0,  8'd34, 9'd292},{1'b0,  8'd47, 9'd182},{1'b0,  8'd72,   9'd0},{1'b0,  8'd73, 9'd169},{1'b0,  8'd97, 9'd175},{1'b0, 8'd117,   9'd0},{1'b1, 8'd118,   9'd6},
{1'b0,  8'd10, 9'd159},{1'b0,  8'd14, 9'd349},{1'b0,  8'd14, 9'd194},{1'b0,  8'd25, 9'd158},{1'b0,  8'd28,   9'd0},{1'b0,  8'd43, 9'd190},{1'b0,  8'd71,  9'd95},{1'b0,  8'd73,   9'd0},{1'b0,  8'd75, 9'd291},{1'b0, 8'd112, 9'd188},{1'b0, 8'd118,   9'd0},{1'b1, 8'd128, 9'd311},
{1'b0,   8'd0,  9'd55},{1'b0,   8'd5, 9'd126},{1'b0,  8'd11,   9'd2},{1'b0,  8'd12,  9'd32},{1'b0,  8'd18,  9'd44},{1'b0,  8'd29,   9'd0},{1'b0,  8'd49,  9'd33},{1'b0,  8'd74,   9'd0},{1'b0,  8'd80,  9'd64},{1'b0,  8'd92, 9'd286},{1'b0, 8'd104, 9'd170},{1'b1, 8'd119,   9'd0},
{1'b0,   8'd3,  9'd34},{1'b0,   8'd6,  9'd75},{1'b0,   8'd6, 9'd132},{1'b0,  8'd10, 9'd165},{1'b0,  8'd20,  9'd87},{1'b0,  8'd30,   9'd0},{1'b0,  8'd65, 9'd313},{1'b0,  8'd70, 9'd123},{1'b0,  8'd75,   9'd0},{1'b0,  8'd91, 9'd307},{1'b0, 8'd120,   9'd0},{1'b1, 8'd126, 9'd143},
{1'b0,   8'd0, 9'd324},{1'b0,   8'd4, 9'd338},{1'b0,   8'd7,  9'd98},{1'b0,  8'd13,  9'd93},{1'b0,  8'd31,   9'd0},{1'b0,  8'd44,  9'd59},{1'b0,  8'd59,  9'd31},{1'b0,  8'd71, 9'd280},{1'b0,  8'd76,   9'd0},{1'b0,  8'd99, 9'd231},{1'b0, 8'd121,   9'd0},{1'b1, 8'd134, 9'd322},
{1'b0,   8'd1, 9'd253},{1'b0,   8'd2, 9'd174},{1'b0,   8'd3,  9'd84},{1'b0,   8'd8,  9'd77},{1'b0,  8'd17, 9'd296},{1'b0,  8'd32,   9'd0},{1'b0,  8'd45,  9'd22},{1'b0,  8'd70, 9'd140},{1'b0,  8'd77,   9'd0},{1'b0, 8'd119, 9'd148},{1'b0, 8'd122,   9'd0},{1'b1, 8'd127, 9'd152},
{1'b0,  8'd10, 9'd225},{1'b0,  8'd14, 9'd248},{1'b0,  8'd14, 9'd335},{1'b0,  8'd33,   9'd0},{1'b0,  8'd37,  9'd45},{1'b0,  8'd42, 9'd138},{1'b0,  8'd52, 9'd269},{1'b0,  8'd65,  9'd28},{1'b0,  8'd78,   9'd0},{1'b0,  8'd95, 9'd204},{1'b0, 8'd123,   9'd0},{1'b1, 8'd130, 9'd107},
{1'b0,   8'd2, 9'd298},{1'b0,   8'd7, 9'd165},{1'b0,  8'd12, 9'd352},{1'b0,  8'd34,   9'd0},{1'b0,  8'd34,  9'd54},{1'b0,  8'd37,  9'd23},{1'b0,  8'd58,  9'd91},{1'b0,  8'd61, 9'd251},{1'b0,  8'd79,   9'd0},{1'b0, 8'd105, 9'd290},{1'b0, 8'd109, 9'd127},{1'b1, 8'd124,   9'd0},
{1'b0,   8'd3, 9'd128},{1'b0,   8'd5,  9'd35},{1'b0,  8'd11,   9'd4},{1'b0,  8'd14, 9'd285},{1'b0,  8'd26, 9'd303},{1'b0,  8'd35,   9'd0},{1'b0,  8'd53, 9'd143},{1'b0,  8'd80,   9'd0},{1'b0,  8'd86, 9'd173},{1'b0, 8'd112, 9'd307},{1'b0, 8'd122, 9'd358},{1'b1, 8'd125,   9'd0},
{1'b0,   8'd3, 9'd174},{1'b0,   8'd5, 9'd352},{1'b0,   8'd6, 9'd340},{1'b0,  8'd13, 9'd184},{1'b0,  8'd28,  9'd54},{1'b0,  8'd36,   9'd0},{1'b0,  8'd66, 9'd307},{1'b0,  8'd79, 9'd164},{1'b0,  8'd81,   9'd0},{1'b0, 8'd117,   9'd8},{1'b0, 8'd124, 9'd322},{1'b1, 8'd126,   9'd0},
{1'b0,   8'd1, 9'd283},{1'b0,   8'd9,  9'd71},{1'b0,  8'd12,  9'd59},{1'b0,  8'd13, 9'd176},{1'b0,  8'd14, 9'd107},{1'b0,  8'd37,   9'd0},{1'b0,  8'd54, 9'd331},{1'b0,  8'd76, 9'd310},{1'b0,  8'd82,   9'd0},{1'b0, 8'd101, 9'd251},{1'b0, 8'd127,   9'd0},{1'b1, 8'd133, 9'd114},
{1'b0,   8'd7, 9'd281},{1'b0,  8'd10,  9'd10},{1'b0,  8'd14, 9'd303},{1'b0,  8'd21, 9'd138},{1'b0,  8'd33, 9'd243},{1'b0,  8'd38,   9'd0},{1'b0,  8'd64,  9'd64},{1'b0,  8'd83,   9'd0},{1'b0,  8'd88, 9'd192},{1'b0, 8'd125, 9'd249},{1'b0, 8'd128,   9'd0},{1'b1, 8'd130, 9'd265},
{1'b0,   8'd0, 9'd163},{1'b0,   8'd7,  9'd46},{1'b0,  8'd10, 9'd291},{1'b0,  8'd19,  9'd95},{1'b0,  8'd32, 9'd133},{1'b0,  8'd39,   9'd0},{1'b0,  8'd49,   9'd7},{1'b0,  8'd83, 9'd107},{1'b0,  8'd84,   9'd0},{1'b0, 8'd101, 9'd205},{1'b0, 8'd111,  9'd29},{1'b1, 8'd129,   9'd0},
{1'b0,   8'd0, 9'd141},{1'b0,   8'd0, 9'd248},{1'b0,  8'd11, 9'd235},{1'b0,  8'd12, 9'd158},{1'b0,  8'd13,  9'd84},{1'b0,  8'd40,   9'd0},{1'b0,  8'd61, 9'd139},{1'b0,  8'd67,  9'd88},{1'b0,  8'd85,   9'd0},{1'b0, 8'd103,  9'd58},{1'b0, 8'd121, 9'd319},{1'b1, 8'd130,   9'd0},
{1'b0,   8'd5, 9'd209},{1'b0,   8'd8, 9'd186},{1'b0,  8'd11, 9'd176},{1'b0,  8'd13,  9'd17},{1'b0,  8'd41,   9'd0},{1'b0,  8'd44, 9'd260},{1'b0,  8'd72, 9'd271},{1'b0,  8'd83, 9'd246},{1'b0,  8'd86,   9'd0},{1'b0,  8'd95, 9'd130},{1'b0, 8'd131,   9'd0},{1'b1, 8'd132, 9'd178},
{1'b0,   8'd1,   9'd7},{1'b0,   8'd1,  9'd18},{1'b0,   8'd3, 9'd194},{1'b0,  8'd24, 9'd314},{1'b0,  8'd24,  9'd65},{1'b0,  8'd42,   9'd0},{1'b0,  8'd54, 9'd281},{1'b0,  8'd63, 9'd201},{1'b0,  8'd87,   9'd0},{1'b0,  8'd93, 9'd181},{1'b0, 8'd117, 9'd109},{1'b1, 8'd132,   9'd0},
{1'b0,   8'd1,  9'd59},{1'b0,   8'd2,  9'd37},{1'b0,   8'd4,  9'd46},{1'b0,  8'd11, 9'd167},{1'b0,  8'd41, 9'd101},{1'b0,  8'd43,   9'd0},{1'b0,  8'd72, 9'd258},{1'b0,  8'd74, 9'd313},{1'b0,  8'd88,   9'd0},{1'b0, 8'd115, 9'd332},{1'b0, 8'd115, 9'd196},{1'b1, 8'd133,   9'd0},
{1'b0,   8'd1, 9'd160},{1'b0,   8'd7,  9'd13},{1'b0,  8'd12, 9'd113},{1'b0,  8'd15,  9'd69},{1'b0,  8'd43, 9'd174},{1'b0,  8'd44,   9'd0},{1'b0,  8'd60, 9'd168},{1'b0,  8'd75, 9'd212},{1'b0,  8'd89,   9'd0},{1'b0,  8'd93,  9'd38},{1'b0, 8'd131, 9'd135},{1'b1, 8'd134,   9'd0}
};
localparam int          cLARGE_HS_TAB_4BY5_PACKED_SIZE = 573;
localparam bit [17 : 0] cLARGE_HS_TAB_4BY5_PACKED[cLARGE_HS_TAB_4BY5_PACKED_SIZE] = '{
{1'b0,   8'd0,   9'd0},{1'b0,   8'd6, 9'd104},{1'b0,  8'd12, 9'd325},{1'b0,  8'd15, 9'd319},{1'b0,  8'd15, 9'd181},{1'b0,  8'd17, 9'd243},{1'b0,  8'd25, 9'd121},{1'b0,  8'd36,   9'd0},{1'b0,  8'd39,  9'd61},{1'b0,  8'd49,  9'd72},{1'b0,  8'd72,   9'd0},{1'b0,  8'd81,  9'd34},{1'b0,  8'd86, 9'd200},{1'b0, 8'd108,   9'd0},{1'b0, 8'd125, 9'd231},{1'b1, 8'd139, 9'd258},
{1'b0,   8'd1,   9'd0},{1'b0,   8'd9,   9'd7},{1'b0,  8'd10, 9'd242},{1'b0,  8'd14,  9'd96},{1'b0,  8'd17, 9'd315},{1'b0,  8'd27, 9'd330},{1'b0,  8'd33, 9'd289},{1'b0,  8'd37,   9'd0},{1'b0,  8'd41, 9'd297},{1'b0,  8'd63,  9'd97},{1'b0,  8'd73,   9'd0},{1'b0,  8'd96,  9'd23},{1'b0,  8'd98, 9'd359},{1'b0, 8'd109,   9'd0},{1'b0, 8'd118, 9'd344},{1'b1, 8'd121, 9'd211},
{1'b0,   8'd2,   9'd0},{1'b0,   8'd5,  9'd95},{1'b0,   8'd7,  9'd31},{1'b0,  8'd10, 9'd218},{1'b0,  8'd12, 9'd107},{1'b0,  8'd19,  9'd28},{1'b0,  8'd21, 9'd341},{1'b0,  8'd38,   9'd0},{1'b0,  8'd48, 9'd332},{1'b0,  8'd67,  9'd58},{1'b0,  8'd74,   9'd0},{1'b0,  8'd78, 9'd156},{1'b0, 8'd106, 9'd226},{1'b0, 8'd110,   9'd0},{1'b0, 8'd118, 9'd333},{1'b1, 8'd125, 9'd183},
{1'b0,   8'd3,   9'd0},{1'b0,   8'd5,  9'd59},{1'b0,   8'd5,  9'd28},{1'b0,   8'd9,  9'd65},{1'b0,  8'd11, 9'd254},{1'b0,  8'd15,  9'd76},{1'b0,  8'd18, 9'd282},{1'b0,  8'd39,   9'd0},{1'b0,  8'd40, 9'd209},{1'b0,  8'd58, 9'd216},{1'b0,  8'd72, 9'd137},{1'b0,  8'd75,   9'd0},{1'b0,  8'd94, 9'd184},{1'b0, 8'd111,   9'd0},{1'b0, 8'd128,   9'd7},{1'b1, 8'd129, 9'd162},
{1'b0,   8'd4,   9'd0},{1'b0,   8'd4, 9'd333},{1'b0,   8'd6,  9'd26},{1'b0,   8'd7, 9'd180},{1'b0,  8'd15, 9'd184},{1'b0,  8'd30,  9'd62},{1'b0,  8'd31, 9'd176},{1'b0,  8'd40,   9'd0},{1'b0,  8'd49, 9'd206},{1'b0,  8'd54, 9'd167},{1'b0,  8'd76,   9'd0},{1'b0,  8'd84,  9'd90},{1'b0, 8'd104,  9'd17},{1'b0, 8'd112,   9'd0},{1'b0, 8'd122,   9'd3},{1'b1, 8'd134, 9'd270},
{1'b0,   8'd0,   9'd4},{1'b0,   8'd5,   9'd0},{1'b0,   8'd5, 9'd113},{1'b0,   8'd9, 9'd125},{1'b0,  8'd13, 9'd318},{1'b0,  8'd16, 9'd229},{1'b0,  8'd22, 9'd122},{1'b0,  8'd41,   9'd0},{1'b0,  8'd44, 9'd223},{1'b0,  8'd51,  9'd19},{1'b0,  8'd77,   9'd0},{1'b0,  8'd97,  9'd61},{1'b0, 8'd105, 9'd271},{1'b0, 8'd113,   9'd0},{1'b0, 8'd128,   9'd3},{1'b1, 8'd129, 9'd172},
{1'b0,   8'd6,   9'd0},{1'b0,   8'd7, 9'd218},{1'b0,   8'd8, 9'd234},{1'b0,  8'd11,  9'd63},{1'b0,  8'd11, 9'd168},{1'b0,  8'd13,  9'd69},{1'b0,  8'd27,  9'd70},{1'b0,  8'd42,   9'd0},{1'b0,  8'd42,  9'd75},{1'b0,  8'd57, 9'd111},{1'b0,  8'd78,   9'd0},{1'b0,  8'd88, 9'd342},{1'b0,  8'd88,  9'd61},{1'b0, 8'd114,   9'd0},{1'b0, 8'd132, 9'd152},{1'b1, 8'd135, 9'd320},
{1'b0,   8'd4, 9'd335},{1'b0,   8'd6,  9'd78},{1'b0,   8'd7,   9'd0},{1'b0,  8'd10, 9'd188},{1'b0,  8'd10, 9'd227},{1'b0,  8'd14, 9'd175},{1'b0,  8'd19, 9'd291},{1'b0,  8'd43,   9'd0},{1'b0,  8'd45, 9'd123},{1'b0,  8'd63,  9'd68},{1'b0,  8'd73, 9'd117},{1'b0,  8'd79,   9'd0},{1'b0,  8'd86,  9'd91},{1'b0, 8'd115,   9'd0},{1'b0, 8'd116, 9'd206},{1'b1, 8'd136, 9'd264},
{1'b0,   8'd0, 9'd225},{1'b0,   8'd8,   9'd0},{1'b0,   8'd8, 9'd262},{1'b0,   8'd9,  9'd43},{1'b0,  8'd10, 9'd248},{1'b0,  8'd14, 9'd105},{1'b0,  8'd20, 9'd247},{1'b0,  8'd44,   9'd0},{1'b0,  8'd52,  9'd36},{1'b0,  8'd70, 9'd236},{1'b0,  8'd77, 9'd249},{1'b0,  8'd80,   9'd0},{1'b0, 8'd100, 9'd165},{1'b0, 8'd112,  9'd96},{1'b0, 8'd116,   9'd0},{1'b1, 8'd133,  9'd59},
{1'b0,   8'd0, 9'd236},{1'b0,   8'd1, 9'd286},{1'b0,   8'd2, 9'd154},{1'b0,   8'd2, 9'd291},{1'b0,   8'd9,   9'd0},{1'b0,  8'd13, 9'd162},{1'b0,  8'd26, 9'd198},{1'b0,  8'd36, 9'd267},{1'b0,  8'd45,   9'd0},{1'b0,  8'd60, 9'd110},{1'b0,  8'd81,   9'd0},{1'b0,  8'd99, 9'd243},{1'b0, 8'd106, 9'd288},{1'b0, 8'd117,   9'd0},{1'b0, 8'd123, 9'd221},{1'b1, 8'd143, 9'd154},
{1'b0,   8'd3,  9'd90},{1'b0,   8'd4, 9'd171},{1'b0,  8'd10,   9'd0},{1'b0,  8'd12, 9'd110},{1'b0,  8'd12,  9'd60},{1'b0,  8'd13, 9'd332},{1'b0,  8'd25, 9'd264},{1'b0,  8'd46,   9'd0},{1'b0,  8'd47, 9'd182},{1'b0,  8'd65, 9'd183},{1'b0,  8'd81, 9'd246},{1'b0,  8'd82,   9'd0},{1'b0,  8'd92, 9'd286},{1'b0, 8'd118,   9'd0},{1'b0, 8'd120, 9'd282},{1'b1, 8'd122,  9'd40},
{1'b0,   8'd8, 9'd114},{1'b0,   8'd8, 9'd238},{1'b0,  8'd11,   9'd0},{1'b0,  8'd12, 9'd358},{1'b0,  8'd15, 9'd336},{1'b0,  8'd15,  9'd15},{1'b0,  8'd33, 9'd324},{1'b0,  8'd47,   9'd0},{1'b0,  8'd56, 9'd123},{1'b0,  8'd65, 9'd319},{1'b0,  8'd75, 9'd151},{1'b0,  8'd83,   9'd0},{1'b0,  8'd90, 9'd266},{1'b0, 8'd119,   9'd0},{1'b0, 8'd126, 9'd250},{1'b1, 8'd136, 9'd342},
{1'b0,   8'd0,  9'd11},{1'b0,   8'd0, 9'd356},{1'b0,   8'd2,  9'd78},{1'b0,  8'd10,  9'd47},{1'b0,  8'd11, 9'd245},{1'b0,  8'd12,   9'd0},{1'b0,  8'd30, 9'd242},{1'b0,  8'd46, 9'd256},{1'b0,  8'd48,   9'd0},{1'b0,  8'd61, 9'd121},{1'b0,  8'd80, 9'd246},{1'b0,  8'd84,   9'd0},{1'b0,  8'd85, 9'd162},{1'b0, 8'd113, 9'd193},{1'b0, 8'd120,   9'd0},{1'b1, 8'd134,  9'd38},
{1'b0,   8'd3,  9'd14},{1'b0,   8'd4, 9'd143},{1'b0,   8'd7, 9'd126},{1'b0,   8'd9, 9'd157},{1'b0,  8'd13,   9'd0},{1'b0,  8'd16,  9'd50},{1'b0,  8'd29, 9'd303},{1'b0,  8'd49,   9'd0},{1'b0,  8'd67, 9'd267},{1'b0,  8'd70,  9'd51},{1'b0,  8'd76,  9'd89},{1'b0,  8'd83, 9'd122},{1'b0,  8'd85,   9'd0},{1'b0, 8'd108, 9'd202},{1'b0, 8'd121,   9'd0},{1'b1, 8'd131,  9'd97},
{1'b0,   8'd7,  9'd35},{1'b0,  8'd11, 9'd331},{1'b0,  8'd14,   9'd0},{1'b0,  8'd15, 9'd226},{1'b0,  8'd17,  9'd58},{1'b0,  8'd22, 9'd196},{1'b0,  8'd32, 9'd238},{1'b0,  8'd50,   9'd0},{1'b0,  8'd62, 9'd148},{1'b0,  8'd69,  9'd99},{1'b0,  8'd83,   9'd7},{1'b0,  8'd86,   9'd0},{1'b0,  8'd87, 9'd313},{1'b0, 8'd122,   9'd0},{1'b0, 8'd127, 9'd261},{1'b1, 8'd130, 9'd358},
{1'b0,   8'd3, 9'd131},{1'b0,   8'd5, 9'd197},{1'b0,   8'd7, 9'd326},{1'b0,   8'd7, 9'd112},{1'b0,  8'd11, 9'd252},{1'b0,  8'd12, 9'd203},{1'b0,  8'd15,   9'd0},{1'b0,  8'd51,   9'd0},{1'b0,  8'd57, 9'd265},{1'b0,  8'd68, 9'd131},{1'b0,  8'd87,   9'd0},{1'b0,  8'd99,  9'd59},{1'b0, 8'd107, 9'd161},{1'b0, 8'd111, 9'd231},{1'b0, 8'd121,  9'd37},{1'b1, 8'd123,   9'd0},
{1'b0,   8'd0, 9'd311},{1'b0,   8'd5, 9'd103},{1'b0,   8'd6, 9'd300},{1'b0,  8'd11, 9'd325},{1'b0,  8'd15,  9'd71},{1'b0,  8'd16,   9'd0},{1'b0,  8'd17, 9'd186},{1'b0,  8'd52,   9'd0},{1'b0,  8'd62, 9'd175},{1'b0,  8'd69,  9'd72},{1'b0,  8'd78, 9'd346},{1'b0,  8'd88,   9'd0},{1'b0, 8'd100, 9'd333},{1'b0, 8'd124,   9'd0},{1'b0, 8'd141,   9'd7},{1'b1, 8'd143, 9'd197},
{1'b0,   8'd1, 9'd145},{1'b0,   8'd1, 9'd107},{1'b0,   8'd6, 9'd321},{1'b0,   8'd8,  9'd11},{1'b0,  8'd17,   9'd0},{1'b0,  8'd17, 9'd152},{1'b0,  8'd46, 9'd115},{1'b0,  8'd53,   9'd0},{1'b0,  8'd68,  9'd64},{1'b0,  8'd79,  9'd40},{1'b0,  8'd89,   9'd0},{1'b0,  8'd96, 9'd269},{1'b0, 8'd124, 9'd248},{1'b0, 8'd124, 9'd205},{1'b1, 8'd125,   9'd0},
{1'b0,   8'd0, 9'd278},{1'b0,   8'd8, 9'd344},{1'b0,   8'd9, 9'd253},{1'b0,  8'd12, 9'd229},{1'b0,  8'd16, 9'd181},{1'b0,  8'd18,   9'd0},{1'b0,  8'd35,  9'd88},{1'b0,  8'd53, 9'd331},{1'b0,  8'd54,   9'd0},{1'b0,  8'd59,  9'd41},{1'b0,  8'd90,   9'd0},{1'b0,  8'd93, 9'd307},{1'b0, 8'd104, 9'd198},{1'b0, 8'd123, 9'd235},{1'b0, 8'd126,   9'd0},{1'b1, 8'd127, 9'd171},
{1'b0,   8'd2, 9'd216},{1'b0,   8'd4,  9'd37},{1'b0,   8'd5, 9'd159},{1'b0,  8'd11, 9'd151},{1'b0,  8'd16, 9'd128},{1'b0,  8'd19,   9'd0},{1'b0,  8'd21, 9'd284},{1'b0,  8'd38, 9'd135},{1'b0,  8'd54, 9'd265},{1'b0,  8'd55,   9'd0},{1'b0,  8'd82, 9'd232},{1'b0,  8'd91,   9'd0},{1'b0,  8'd97,  9'd50},{1'b0, 8'd110, 9'd250},{1'b0, 8'd119, 9'd270},{1'b1, 8'd127,   9'd0},
{1'b0,   8'd2, 9'd336},{1'b0,   8'd2,  9'd82},{1'b0,   8'd3, 9'd119},{1'b0,  8'd14, 9'd221},{1'b0,  8'd17,  9'd81},{1'b0,  8'd20,   9'd0},{1'b0,  8'd29,  9'd84},{1'b0,  8'd39,   9'd9},{1'b0,  8'd52,  9'd25},{1'b0,  8'd56,   9'd0},{1'b0,  8'd79,  9'd35},{1'b0,  8'd92,   9'd0},{1'b0, 8'd107, 9'd211},{1'b0, 8'd117, 9'd225},{1'b0, 8'd128,   9'd0},{1'b1, 8'd139,  9'd85},
{1'b0,   8'd1, 9'd296},{1'b0,  8'd13, 9'd311},{1'b0,  8'd14, 9'd214},{1'b0,  8'd14, 9'd166},{1'b0,  8'd17, 9'd345},{1'b0,  8'd21,   9'd0},{1'b0,  8'd26, 9'd285},{1'b0,  8'd56, 9'd116},{1'b0,  8'd57,   9'd0},{1'b0,  8'd60, 9'd298},{1'b0,  8'd77,  9'd18},{1'b0,  8'd92, 9'd334},{1'b0,  8'd93,   9'd0},{1'b0, 8'd116, 9'd155},{1'b0, 8'd129,   9'd0},{1'b1, 8'd131, 9'd121},
{1'b0,   8'd1,  9'd13},{1'b0,   8'd6, 9'd264},{1'b0,   8'd6, 9'd319},{1'b0,  8'd16, 9'd168},{1'b0,  8'd16, 9'd103},{1'b0,  8'd22,   9'd0},{1'b0,  8'd43, 9'd166},{1'b0,  8'd45, 9'd134},{1'b0,  8'd58,   9'd0},{1'b0,  8'd75, 9'd193},{1'b0,  8'd76, 9'd156},{1'b0,  8'd94,   9'd0},{1'b0, 8'd111, 9'd122},{1'b0, 8'd130,   9'd0},{1'b1, 8'd138, 9'd250},
{1'b0,   8'd4, 9'd338},{1'b0,   8'd4,  9'd65},{1'b0,   8'd7, 9'd319},{1'b0,   8'd7, 9'd144},{1'b0,  8'd23,   9'd0},{1'b0,  8'd34, 9'd179},{1'b0,  8'd42, 9'd187},{1'b0,  8'd59,   9'd0},{1'b0,  8'd61,  9'd96},{1'b0,  8'd89, 9'd125},{1'b0,  8'd95,   9'd0},{1'b0, 8'd101,  9'd88},{1'b0, 8'd113,  9'd56},{1'b0, 8'd131,   9'd0},{1'b1, 8'd137, 9'd228},
{1'b0,   8'd0, 9'd176},{1'b0,   8'd2,  9'd15},{1'b0,   8'd5, 9'd189},{1'b0,   8'd5, 9'd306},{1'b0,  8'd11, 9'd120},{1'b0,  8'd15, 9'd273},{1'b0,  8'd24,   9'd0},{1'b0,  8'd50, 9'd267},{1'b0,  8'd55,   9'd8},{1'b0,  8'd60,   9'd0},{1'b0,  8'd74, 9'd304},{1'b0,  8'd96,   9'd0},{1'b0, 8'd103, 9'd197},{1'b0, 8'd109, 9'd215},{1'b0, 8'd132,   9'd0},{1'b1, 8'd137,  9'd48},
{1'b0,   8'd3, 9'd280},{1'b0,  8'd13,  9'd22},{1'b0,  8'd14, 9'd125},{1'b0,  8'd17, 9'd217},{1'b0,  8'd17, 9'd332},{1'b0,  8'd25,   9'd0},{1'b0,  8'd28,  9'd54},{1'b0,  8'd61,   9'd0},{1'b0,  8'd64, 9'd337},{1'b0,  8'd64, 9'd205},{1'b0,  8'd95, 9'd274},{1'b0,  8'd97,   9'd0},{1'b0, 8'd102, 9'd303},{1'b0, 8'd117, 9'd135},{1'b0, 8'd133,   9'd0},{1'b1, 8'd133, 9'd123},
{1'b0,   8'd1, 9'd103},{1'b0,   8'd6,  9'd40},{1'b0,   8'd9, 9'd115},{1'b0,  8'd10, 9'd228},{1'b0,  8'd13, 9'd122},{1'b0,  8'd20, 9'd284},{1'b0,  8'd26,   9'd0},{1'b0,  8'd40, 9'd184},{1'b0,  8'd50, 9'd244},{1'b0,  8'd62,   9'd0},{1'b0,  8'd74, 9'd223},{1'b0,  8'd87,  9'd41},{1'b0,  8'd98,   9'd0},{1'b0, 8'd115,  9'd19},{1'b0, 8'd119, 9'd278},{1'b1, 8'd134,   9'd0},
{1'b0,   8'd6, 9'd312},{1'b0,   8'd8, 9'd123},{1'b0,   8'd9, 9'd130},{1'b0,  8'd10, 9'd246},{1'b0,  8'd13,  9'd40},{1'b0,  8'd15, 9'd111},{1'b0,  8'd27,   9'd0},{1'b0,  8'd44, 9'd306},{1'b0,  8'd63,   9'd0},{1'b0,  8'd66, 9'd123},{1'b0,  8'd85, 9'd167},{1'b0,  8'd90, 9'd194},{1'b0,  8'd99,   9'd0},{1'b0, 8'd135,   9'd0},{1'b0, 8'd140, 9'd208},{1'b1, 8'd142, 9'd111},
{1'b0,   8'd3,  9'd19},{1'b0,   8'd3, 9'd208},{1'b0,   8'd5, 9'd298},{1'b0,   8'd6,  9'd33},{1'b0,  8'd17, 9'd212},{1'b0,  8'd24, 9'd332},{1'b0,  8'd28,   9'd0},{1'b0,  8'd41,  9'd67},{1'b0,  8'd58, 9'd339},{1'b0,  8'd64,   9'd0},{1'b0,  8'd93, 9'd141},{1'b0, 8'd100,   9'd0},{1'b0, 8'd101, 9'd241},{1'b0, 8'd120,  9'd11},{1'b0, 8'd130, 9'd106},{1'b1, 8'd136,   9'd0},
{1'b0,   8'd2, 9'd196},{1'b0,  8'd12, 9'd263},{1'b0,  8'd13,  9'd14},{1'b0,  8'd14,  9'd42},{1'b0,  8'd16, 9'd219},{1'b0,  8'd28, 9'd318},{1'b0,  8'd29,   9'd0},{1'b0,  8'd53,  9'd34},{1'b0,  8'd55, 9'd210},{1'b0,  8'd65,   9'd0},{1'b0,  8'd89,  9'd26},{1'b0,  8'd98, 9'd185},{1'b0, 8'd101,   9'd0},{1'b0, 8'd137,   9'd0},{1'b0, 8'd138,  9'd13},{1'b1, 8'd142, 9'd342},
{1'b0,   8'd1, 9'd138},{1'b0,   8'd2, 9'd242},{1'b0,   8'd8,  9'd62},{1'b0,  8'd14,  9'd82},{1'b0,  8'd16, 9'd341},{1'b0,  8'd30,   9'd0},{1'b0,  8'd35, 9'd338},{1'b0,  8'd47, 9'd340},{1'b0,  8'd51, 9'd150},{1'b0,  8'd66,   9'd0},{1'b0,  8'd94, 9'd191},{1'b0, 8'd102,   9'd0},{1'b0, 8'd105, 9'd142},{1'b0, 8'd112,  9'd17},{1'b0, 8'd114,  9'd21},{1'b1, 8'd138,   9'd0},
{1'b0,   8'd0, 9'd154},{1'b0,   8'd0, 9'd348},{1'b0,   8'd8, 9'd219},{1'b0,  8'd13, 9'd145},{1'b0,  8'd23, 9'd340},{1'b0,  8'd31,   9'd0},{1'b0,  8'd34, 9'd354},{1'b0,  8'd37, 9'd155},{1'b0,  8'd67,   9'd0},{1'b0,  8'd71, 9'd111},{1'b0,  8'd72, 9'd156},{1'b0,  8'd80, 9'd107},{1'b0, 8'd103,   9'd0},{1'b0, 8'd109, 9'd301},{1'b0, 8'd110, 9'd342},{1'b1, 8'd139,   9'd0},
{1'b0,   8'd1,  9'd85},{1'b0,   8'd8, 9'd195},{1'b0,  8'd11, 9'd312},{1'b0,  8'd14, 9'd264},{1'b0,  8'd24, 9'd189},{1'b0,  8'd31, 9'd252},{1'b0,  8'd32,   9'd0},{1'b0,  8'd43, 9'd142},{1'b0,  8'd48, 9'd210},{1'b0,  8'd68,   9'd0},{1'b0,  8'd82, 9'd165},{1'b0,  8'd91,  9'd70},{1'b0, 8'd104,   9'd0},{1'b0, 8'd132, 9'd240},{1'b0, 8'd140,   9'd0},{1'b1, 8'd141,  9'd74},
{1'b0,   8'd2,  9'd59},{1'b0,   8'd3,  9'd78},{1'b0,   8'd4,  9'd14},{1'b0,   8'd9, 9'd107},{1'b0,  8'd12, 9'd286},{1'b0,  8'd16,  9'd48},{1'b0,  8'd33,   9'd0},{1'b0,  8'd36, 9'd317},{1'b0,  8'd66, 9'd327},{1'b0,  8'd69,   9'd0},{1'b0,  8'd95,  9'd58},{1'b0, 8'd103, 9'd174},{1'b0, 8'd105,   9'd0},{1'b0, 8'd114,  9'd83},{1'b0, 8'd140,  9'd68},{1'b1, 8'd141,   9'd0},
{1'b0,   8'd3, 9'd231},{1'b0,   8'd4, 9'd117},{1'b0,   8'd9, 9'd103},{1'b0,  8'd10, 9'd220},{1'b0,  8'd18, 9'd116},{1'b0,  8'd32, 9'd203},{1'b0,  8'd34,   9'd0},{1'b0,  8'd37, 9'd207},{1'b0,  8'd59, 9'd243},{1'b0,  8'd70,   9'd0},{1'b0,  8'd73,  9'd51},{1'b0,  8'd84, 9'd102},{1'b0, 8'd106,   9'd0},{1'b0, 8'd115,  9'd57},{1'b0, 8'd126, 9'd189},{1'b1, 8'd142,   9'd0},
{1'b0,   8'd1, 9'd213},{1'b0,   8'd3,  9'd74},{1'b0,   8'd4, 9'd312},{1'b0,  8'd10, 9'd239},{1'b0,  8'd12,  9'd57},{1'b0,  8'd23, 9'd107},{1'b0,  8'd35,   9'd0},{1'b0,  8'd38, 9'd119},{1'b0,  8'd71,   9'd0},{1'b0,  8'd71,  9'd31},{1'b0,  8'd91,  9'd56},{1'b0, 8'd102, 9'd226},{1'b0, 8'd107,   9'd0},{1'b0, 8'd108, 9'd273},{1'b0, 8'd135, 9'd336},{1'b1, 8'd143,   9'd0}
};
localparam int          cLARGE_HS_TAB_5BY6_PACKED_SIZE = 590;
localparam bit [17 : 0] cLARGE_HS_TAB_5BY6_PACKED[cLARGE_HS_TAB_5BY6_PACKED_SIZE] = '{
{1'b0,   8'd0,   9'd0},{1'b0,   8'd3, 9'd312},{1'b0,   8'd6, 9'd332},{1'b0,   8'd8,  9'd86},{1'b0,   8'd9, 9'd128},{1'b0,  8'd13, 9'd142},{1'b0,  8'd14, 9'd120},{1'b0,  8'd14,  9'd19},{1'b0,  8'd30,   9'd0},{1'b0,  8'd40,  9'd88},{1'b0,  8'd54, 9'd280},{1'b0,  8'd60,   9'd0},{1'b0,  8'd72, 9'd280},{1'b0,  8'd78,  9'd21},{1'b0,  8'd90,   9'd0},{1'b0,  8'd97, 9'd108},{1'b0, 8'd118, 9'd161},{1'b0, 8'd120,   9'd0},{1'b0, 8'd136, 9'd111},{1'b1, 8'd140, 9'd151},
{1'b0,   8'd1,   9'd0},{1'b0,   8'd1, 9'd201},{1'b0,   8'd2, 9'd103},{1'b0,   8'd2, 9'd189},{1'b0,   8'd7, 9'd263},{1'b0,  8'd13, 9'd223},{1'b0,  8'd15, 9'd254},{1'b0,  8'd19, 9'd284},{1'b0,  8'd31,   9'd0},{1'b0,  8'd31,  9'd88},{1'b0,  8'd46, 9'd273},{1'b0,  8'd61,   9'd0},{1'b0,  8'd67, 9'd171},{1'b0,  8'd69, 9'd211},{1'b0,  8'd91,   9'd0},{1'b0, 8'd100, 9'd191},{1'b0, 8'd101, 9'd204},{1'b0, 8'd121,   9'd0},{1'b1, 8'd131,  9'd43},
{1'b0,   8'd0,  9'd97},{1'b0,   8'd2,   9'd0},{1'b0,   8'd5, 9'd135},{1'b0,   8'd9, 9'd219},{1'b0,  8'd12, 9'd318},{1'b0,  8'd12, 9'd245},{1'b0,  8'd27, 9'd169},{1'b0,  8'd28, 9'd118},{1'b0,  8'd32,   9'd0},{1'b0,  8'd42, 9'd186},{1'b0,  8'd56, 9'd168},{1'b0,  8'd62,   9'd0},{1'b0,  8'd65, 9'd155},{1'b0,  8'd70, 9'd222},{1'b0,  8'd91, 9'd120},{1'b0,  8'd92,   9'd0},{1'b0, 8'd116,  9'd12},{1'b0, 8'd122,   9'd0},{1'b0, 8'd130, 9'd204},{1'b1, 8'd132, 9'd353},
{1'b0,   8'd0, 9'd224},{1'b0,   8'd3,   9'd0},{1'b0,   8'd4, 9'd328},{1'b0,   8'd5, 9'd123},{1'b0,   8'd8,  9'd96},{1'b0,  8'd11, 9'd353},{1'b0,  8'd12, 9'd354},{1'b0,  8'd17, 9'd243},{1'b0,  8'd33,   9'd0},{1'b0,  8'd34, 9'd250},{1'b0,  8'd58, 9'd240},{1'b0,  8'd63,   9'd0},{1'b0,  8'd64, 9'd217},{1'b0,  8'd79,  9'd12},{1'b0,  8'd90, 9'd105},{1'b0,  8'd93,   9'd0},{1'b0, 8'd111,  9'd25},{1'b0, 8'd123,   9'd0},{1'b1, 8'd137, 9'd352},
{1'b0,   8'd4,   9'd0},{1'b0,   8'd4, 9'd261},{1'b0,   8'd5, 9'd238},{1'b0,   8'd8,  9'd34},{1'b0,   8'd9,  9'd69},{1'b0,   8'd9, 9'd103},{1'b0,  8'd11,  9'd13},{1'b0,  8'd15, 9'd210},{1'b0,  8'd34,   9'd0},{1'b0,  8'd39, 9'd132},{1'b0,  8'd55,  9'd13},{1'b0,  8'd64,   9'd0},{1'b0,  8'd77,  9'd95},{1'b0,  8'd87, 9'd202},{1'b0,  8'd94,   9'd0},{1'b0, 8'd109, 9'd302},{1'b0, 8'd113,  9'd87},{1'b0, 8'd124,   9'd0},{1'b0, 8'd137, 9'd142},{1'b1, 8'd146, 9'd214},
{1'b0,   8'd2, 9'd339},{1'b0,   8'd2, 9'd166},{1'b0,   8'd4, 9'd161},{1'b0,   8'd5,   9'd0},{1'b0,   8'd7, 9'd158},{1'b0,   8'd8,  9'd73},{1'b0,  8'd12,  9'd24},{1'b0,  8'd13, 9'd125},{1'b0,  8'd35,   9'd0},{1'b0,  8'd48, 9'd110},{1'b0,  8'd55, 9'd275},{1'b0,  8'd63, 9'd353},{1'b0,  8'd65,   9'd0},{1'b0,  8'd89,  9'd96},{1'b0,  8'd91, 9'd135},{1'b0,  8'd95,   9'd0},{1'b0, 8'd115,  9'd69},{1'b0, 8'd125,   9'd0},{1'b0, 8'd132, 9'd298},{1'b1, 8'd147, 9'd125},
{1'b0,   8'd0, 9'd107},{1'b0,   8'd3, 9'd333},{1'b0,   8'd6,   9'd0},{1'b0,   8'd6, 9'd277},{1'b0,   8'd7, 9'd139},{1'b0,   8'd9, 9'd126},{1'b0,  8'd11, 9'd121},{1'b0,  8'd17, 9'd226},{1'b0,  8'd36,   9'd0},{1'b0,  8'd37, 9'd309},{1'b0,  8'd45, 9'd150},{1'b0,  8'd66,   9'd0},{1'b0,  8'd73, 9'd305},{1'b0,  8'd86, 9'd151},{1'b0,  8'd96,   9'd0},{1'b0, 8'd107, 9'd267},{1'b0, 8'd111, 9'd244},{1'b0, 8'd126,   9'd0},{1'b0, 8'd129, 9'd322},{1'b1, 8'd143,  9'd70},
{1'b0,   8'd1, 9'd213},{1'b0,   8'd2, 9'd242},{1'b0,   8'd3, 9'd143},{1'b0,   8'd7,   9'd0},{1'b0,   8'd7,  9'd57},{1'b0,  8'd22, 9'd317},{1'b0,  8'd27,  9'd35},{1'b0,  8'd37,   9'd0},{1'b0,  8'd47, 9'd205},{1'b0,  8'd52,  9'd37},{1'b0,  8'd62,   9'd2},{1'b0,  8'd67,   9'd0},{1'b0,  8'd83, 9'd192},{1'b0,  8'd92,  9'd57},{1'b0,  8'd97,   9'd0},{1'b0, 8'd116, 9'd156},{1'b0, 8'd120, 9'd261},{1'b0, 8'd123, 9'd122},{1'b1, 8'd127,   9'd0},
{1'b0,   8'd1, 9'd299},{1'b0,   8'd3, 9'd335},{1'b0,   8'd3, 9'd171},{1'b0,   8'd8,   9'd0},{1'b0,  8'd12, 9'd252},{1'b0,  8'd13, 9'd293},{1'b0,  8'd22, 9'd342},{1'b0,  8'd28, 9'd264},{1'b0,  8'd38,   9'd0},{1'b0,  8'd39,  9'd11},{1'b0,  8'd56, 9'd211},{1'b0,  8'd62, 9'd241},{1'b0,  8'd68,   9'd0},{1'b0,  8'd71, 9'd341},{1'b0,  8'd94, 9'd263},{1'b0,  8'd98,   9'd0},{1'b0, 8'd100, 9'd262},{1'b0, 8'd128,   9'd0},{1'b0, 8'd130, 9'd236},{1'b1, 8'd141, 9'd227},
{1'b0,   8'd2, 9'd300},{1'b0,   8'd4,  9'd79},{1'b0,   8'd6, 9'd173},{1'b0,   8'd6,  9'd23},{1'b0,   8'd8,  9'd56},{1'b0,   8'd8, 9'd148},{1'b0,   8'd9,   9'd0},{1'b0,  8'd13, 9'd247},{1'b0,  8'd39,   9'd0},{1'b0,  8'd53, 9'd187},{1'b0,  8'd58,  9'd66},{1'b0,  8'd69,   9'd0},{1'b0,  8'd77, 9'd282},{1'b0,  8'd82, 9'd302},{1'b0,  8'd98, 9'd316},{1'b0,  8'd99,   9'd0},{1'b0, 8'd105, 9'd100},{1'b0, 8'd121,  9'd56},{1'b0, 8'd129,   9'd0},{1'b1, 8'd133, 9'd120},
{1'b0,   8'd0,  9'd85},{1'b0,   8'd3, 9'd112},{1'b0,   8'd4, 9'd102},{1'b0,   8'd9,  9'd48},{1'b0,  8'd10,   9'd0},{1'b0,  8'd14, 9'd217},{1'b0,  8'd18, 9'd198},{1'b0,  8'd24, 9'd185},{1'b0,  8'd34, 9'd313},{1'b0,  8'd40,   9'd0},{1'b0,  8'd49,  9'd51},{1'b0,  8'd70,   9'd0},{1'b0,  8'd76,  9'd56},{1'b0,  8'd83, 9'd135},{1'b0, 8'd100,   9'd0},{1'b0, 8'd103,  9'd19},{1'b0, 8'd117, 9'd331},{1'b0, 8'd128, 9'd110},{1'b0, 8'd130,   9'd0},{1'b1, 8'd133, 9'd237},
{1'b0,   8'd1, 9'd100},{1'b0,   8'd5, 9'd262},{1'b0,   8'd6, 9'd344},{1'b0,   8'd6,  9'd66},{1'b0,  8'd11,   9'd0},{1'b0,  8'd11, 9'd285},{1'b0,  8'd12,  9'd84},{1'b0,  8'd13, 9'd238},{1'b0,  8'd41,   9'd0},{1'b0,  8'd45, 9'd116},{1'b0,  8'd59,  9'd59},{1'b0,  8'd63, 9'd294},{1'b0,  8'd71,   9'd0},{1'b0,  8'd89,  9'd68},{1'b0,  8'd90, 9'd356},{1'b0, 8'd101,   9'd0},{1'b0, 8'd115,  9'd20},{1'b0, 8'd131,   9'd0},{1'b0, 8'd144, 9'd229},{1'b1, 8'd145,  9'd72},
{1'b0,   8'd0, 9'd145},{1'b0,   8'd2, 9'd136},{1'b0,   8'd7, 9'd358},{1'b0,   8'd9,  9'd50},{1'b0,  8'd10, 9'd315},{1'b0,  8'd11, 9'd129},{1'b0,  8'd12,   9'd0},{1'b0,  8'd29, 9'd125},{1'b0,  8'd37,  9'd56},{1'b0,  8'd42,   9'd0},{1'b0,  8'd46, 9'd139},{1'b0,  8'd72,   9'd0},{1'b0,  8'd81, 9'd223},{1'b0,  8'd86, 9'd296},{1'b0,  8'd98, 9'd222},{1'b0, 8'd102,   9'd0},{1'b0, 8'd102, 9'd304},{1'b0, 8'd132,   9'd0},{1'b0, 8'd135, 9'd268},{1'b1, 8'd146, 9'd135},
{1'b0,   8'd0, 9'd286},{1'b0,   8'd1, 9'd310},{1'b0,   8'd4, 9'd278},{1'b0,   8'd7, 9'd229},{1'b0,   8'd9, 9'd286},{1'b0,  8'd12,  9'd54},{1'b0,  8'd13,   9'd0},{1'b0,  8'd13, 9'd275},{1'b0,  8'd42, 9'd189},{1'b0,  8'd43,   9'd0},{1'b0,  8'd43, 9'd317},{1'b0,  8'd73,   9'd0},{1'b0,  8'd87,  9'd28},{1'b0,  8'd88, 9'd196},{1'b0, 8'd102, 9'd161},{1'b0, 8'd103,   9'd0},{1'b0, 8'd119,  9'd45},{1'b0, 8'd133,   9'd0},{1'b0, 8'd142, 9'd113},{1'b1, 8'd144, 9'd129},
{1'b0,   8'd3,  9'd14},{1'b0,   8'd5,  9'd69},{1'b0,   8'd6,  9'd43},{1'b0,   8'd7, 9'd325},{1'b0,   8'd9, 9'd181},{1'b0,  8'd11, 9'd273},{1'b0,  8'd12,   9'd2},{1'b0,  8'd14,   9'd0},{1'b0,  8'd32,  9'd92},{1'b0,  8'd44,   9'd0},{1'b0,  8'd59, 9'd172},{1'b0,  8'd61, 9'd140},{1'b0,  8'd71, 9'd320},{1'b0,  8'd74,   9'd0},{1'b0, 8'd104,   9'd0},{1'b0, 8'd113, 9'd261},{1'b0, 8'd117, 9'd289},{1'b0, 8'd125, 9'd141},{1'b0, 8'd127, 9'd131},{1'b1, 8'd134,   9'd0},
{1'b0,   8'd0, 9'd213},{1'b0,   8'd5, 9'd114},{1'b0,   8'd5, 9'd219},{1'b0,  8'd10, 9'd332},{1'b0,  8'd11, 9'd264},{1'b0,  8'd14,  9'd66},{1'b0,  8'd15,   9'd0},{1'b0,  8'd25,  9'd18},{1'b0,  8'd31, 9'd321},{1'b0,  8'd45,   9'd0},{1'b0,  8'd51, 9'd222},{1'b0,  8'd72, 9'd267},{1'b0,  8'd75,   9'd0},{1'b0,  8'd80, 9'd137},{1'b0, 8'd105,   9'd0},{1'b0, 8'd106,   9'd6},{1'b0, 8'd108, 9'd306},{1'b0, 8'd126, 9'd341},{1'b0, 8'd135,   9'd0},{1'b1, 8'd136,  9'd96},
{1'b0,   8'd0, 9'd138},{1'b0,   8'd1,  9'd59},{1'b0,   8'd2, 9'd290},{1'b0,   8'd5,  9'd62},{1'b0,   8'd8, 9'd216},{1'b0,  8'd14, 9'd181},{1'b0,  8'd16,   9'd0},{1'b0,  8'd29, 9'd107},{1'b0,  8'd36, 9'd348},{1'b0,  8'd43,  9'd30},{1'b0,  8'd46,   9'd0},{1'b0,  8'd61, 9'd112},{1'b0,  8'd76,   9'd0},{1'b0,  8'd82, 9'd307},{1'b0, 8'd106,   9'd0},{1'b0, 8'd108,  9'd50},{1'b0, 8'd114,  9'd21},{1'b0, 8'd129, 9'd211},{1'b0, 8'd136,   9'd0},{1'b1, 8'd138, 9'd216},
{1'b0,   8'd1,  9'd98},{1'b0,   8'd1, 9'd340},{1'b0,   8'd2,  9'd92},{1'b0,   8'd4,  9'd77},{1'b0,   8'd6, 9'd130},{1'b0,   8'd9, 9'd168},{1'b0,  8'd17,   9'd0},{1'b0,  8'd26, 9'd127},{1'b0,  8'd38, 9'd334},{1'b0,  8'd40, 9'd169},{1'b0,  8'd47,   9'd0},{1'b0,  8'd69, 9'd183},{1'b0,  8'd74, 9'd235},{1'b0,  8'd77,   9'd0},{1'b0,  8'd95,  9'd20},{1'b0,  8'd99, 9'd248},{1'b0, 8'd107,   9'd0},{1'b0, 8'd137,   9'd0},{1'b1, 8'd139, 9'd293},
{1'b0,   8'd3,  9'd37},{1'b0,   8'd5,  9'd11},{1'b0,   8'd7, 9'd129},{1'b0,  8'd10,  9'd61},{1'b0,  8'd11, 9'd332},{1'b0,  8'd14,  9'd25},{1'b0,  8'd16, 9'd216},{1'b0,  8'd18,   9'd0},{1'b0,  8'd38, 9'd134},{1'b0,  8'd41,  9'd28},{1'b0,  8'd48,   9'd0},{1'b0,  8'd67, 9'd262},{1'b0,  8'd78,   9'd0},{1'b0,  8'd80, 9'd233},{1'b0, 8'd105,  9'd75},{1'b0, 8'd108,   9'd0},{1'b0, 8'd119, 9'd234},{1'b0, 8'd123, 9'd330},{1'b0, 8'd134, 9'd305},{1'b1, 8'd138,   9'd0},
{1'b0,   8'd0, 9'd165},{1'b0,   8'd1,  9'd82},{1'b0,   8'd1, 9'd144},{1'b0,   8'd2, 9'd329},{1'b0,   8'd7, 9'd333},{1'b0,  8'd10, 9'd212},{1'b0,  8'd19,   9'd0},{1'b0,  8'd23, 9'd311},{1'b0,  8'd49,   9'd0},{1'b0,  8'd51, 9'd135},{1'b0,  8'd57, 9'd170},{1'b0,  8'd60, 9'd118},{1'b0,  8'd66,  9'd47},{1'b0,  8'd79,   9'd0},{1'b0,  8'd94,  9'd64},{1'b0, 8'd106,  9'd80},{1'b0, 8'd109,   9'd0},{1'b0, 8'd122,  9'd78},{1'b0, 8'd139,   9'd0},{1'b1, 8'd140,  9'd66},
{1'b0,   8'd5, 9'd344},{1'b0,   8'd5, 9'd195},{1'b0,   8'd8, 9'd180},{1'b0,  8'd14,   9'd6},{1'b0,  8'd20,   9'd0},{1'b0,  8'd21,  9'd39},{1'b0,  8'd26, 9'd286},{1'b0,  8'd30,  9'd80},{1'b0,  8'd35,  9'd61},{1'b0,  8'd50,   9'd0},{1'b0,  8'd65, 9'd176},{1'b0,  8'd73, 9'd187},{1'b0,  8'd80,   9'd0},{1'b0,  8'd99, 9'd105},{1'b0, 8'd104, 9'd309},{1'b0, 8'd110,   9'd0},{1'b0, 8'd122, 9'd335},{1'b0, 8'd124, 9'd230},{1'b1, 8'd140,   9'd0},
{1'b0,   8'd4, 9'd243},{1'b0,   8'd6, 9'd103},{1'b0,   8'd6,  9'd53},{1'b0,   8'd8,   9'd3},{1'b0,   8'd9, 9'd110},{1'b0,  8'd14, 9'd225},{1'b0,  8'd21,   9'd0},{1'b0,  8'd23,  9'd72},{1'b0,  8'd33, 9'd177},{1'b0,  8'd33,  9'd67},{1'b0,  8'd51,   9'd0},{1'b0,  8'd64,  9'd40},{1'b0,  8'd70, 9'd164},{1'b0,  8'd81,   9'd0},{1'b0, 8'd103, 9'd319},{1'b0, 8'd111,   9'd0},{1'b0, 8'd112, 9'd209},{1'b0, 8'd121, 9'd126},{1'b0, 8'd126, 9'd260},{1'b1, 8'd141,   9'd0},
{1'b0,   8'd0, 9'd103},{1'b0,   8'd3, 9'd301},{1'b0,   8'd9, 9'd329},{1'b0,  8'd10, 9'd345},{1'b0,  8'd13,  9'd82},{1'b0,  8'd13,  9'd69},{1'b0,  8'd14, 9'd296},{1'b0,  8'd22,   9'd0},{1'b0,  8'd32,  9'd81},{1'b0,  8'd47, 9'd339},{1'b0,  8'd52,   9'd0},{1'b0,  8'd81,  9'd53},{1'b0,  8'd82,   9'd0},{1'b0,  8'd85, 9'd185},{1'b0, 8'd101, 9'd357},{1'b0, 8'd109, 9'd268},{1'b0, 8'd112,   9'd0},{1'b0, 8'd134, 9'd303},{1'b0, 8'd141, 9'd306},{1'b1, 8'd142,   9'd0},
{1'b0,   8'd8, 9'd200},{1'b0,  8'd10, 9'd243},{1'b0,  8'd13, 9'd166},{1'b0,  8'd13, 9'd306},{1'b0,  8'd14,  9'd36},{1'b0,  8'd19,  9'd59},{1'b0,  8'd21, 9'd325},{1'b0,  8'd23,   9'd0},{1'b0,  8'd41, 9'd115},{1'b0,  8'd53,   9'd0},{1'b0,  8'd54, 9'd282},{1'b0,  8'd79, 9'd181},{1'b0,  8'd83,   9'd0},{1'b0,  8'd84, 9'd124},{1'b0, 8'd112, 9'd127},{1'b0, 8'd113,   9'd0},{1'b0, 8'd114,  9'd76},{1'b0, 8'd135, 9'd206},{1'b0, 8'd143,   9'd0},{1'b1, 8'd143, 9'd300},
{1'b0,   8'd1, 9'd182},{1'b0,   8'd2, 9'd295},{1'b0,   8'd3, 9'd130},{1'b0,   8'd4,  9'd26},{1'b0,   8'd7, 9'd153},{1'b0,  8'd20, 9'd205},{1'b0,  8'd20, 9'd261},{1'b0,  8'd24,   9'd0},{1'b0,  8'd36, 9'd325},{1'b0,  8'd54,   9'd0},{1'b0,  8'd57, 9'd205},{1'b0,  8'd60,  9'd48},{1'b0,  8'd68, 9'd342},{1'b0,  8'd84,   9'd0},{1'b0,  8'd96, 9'd284},{1'b0,  8'd96,  9'd45},{1'b0, 8'd114,   9'd0},{1'b0, 8'd124,  9'd63},{1'b0, 8'd142,  9'd57},{1'b1, 8'd144,   9'd0},
{1'b0,   8'd3, 9'd159},{1'b0,   8'd3, 9'd338},{1'b0,  8'd10, 9'd152},{1'b0,  8'd11,  9'd79},{1'b0,  8'd12, 9'd259},{1'b0,  8'd12, 9'd303},{1'b0,  8'd13, 9'd336},{1'b0,  8'd25,   9'd0},{1'b0,  8'd30, 9'd234},{1'b0,  8'd53, 9'd102},{1'b0,  8'd55,   9'd0},{1'b0,  8'd68, 9'd147},{1'b0,  8'd75, 9'd113},{1'b0,  8'd85,   9'd0},{1'b0, 8'd110,  9'd69},{1'b0, 8'd115,   9'd0},{1'b0, 8'd118,  9'd68},{1'b0, 8'd139, 9'd254},{1'b0, 8'd145,   9'd0},{1'b1, 8'd145, 9'd129},
{1'b0,   8'd0,  9'd13},{1'b0,   8'd6, 9'd115},{1'b0,  8'd10, 9'd217},{1'b0,  8'd10,  9'd58},{1'b0,  8'd25,  9'd51},{1'b0,  8'd26,   9'd0},{1'b0,  8'd50, 9'd158},{1'b0,  8'd52,  9'd33},{1'b0,  8'd56,   9'd0},{1'b0,  8'd76, 9'd128},{1'b0,  8'd78, 9'd206},{1'b0,  8'd86,   9'd0},{1'b0,  8'd95,   9'd6},{1'b0,  8'd97, 9'd355},{1'b0, 8'd116,   9'd0},{1'b0, 8'd138, 9'd351},{1'b0, 8'd146,   9'd0},{1'b1, 8'd147, 9'd317},
{1'b0,   8'd4, 9'd238},{1'b0,   8'd7, 9'd107},{1'b0,   8'd8, 9'd352},{1'b0,  8'd11, 9'd308},{1'b0,  8'd12, 9'd228},{1'b0,  8'd12, 9'd213},{1'b0,  8'd14, 9'd150},{1'b0,  8'd27,   9'd0},{1'b0,  8'd44, 9'd136},{1'b0,  8'd50,  9'd89},{1'b0,  8'd57,   9'd0},{1'b0,  8'd75, 9'd300},{1'b0,  8'd84, 9'd307},{1'b0,  8'd87,   9'd0},{1'b0, 8'd104, 9'd208},{1'b0, 8'd107,  9'd51},{1'b0, 8'd117,   9'd0},{1'b0, 8'd131, 9'd260},{1'b1, 8'd147,   9'd0},
{1'b0,   8'd1, 9'd242},{1'b0,   8'd4,  9'd50},{1'b0,   8'd8,  9'd98},{1'b0,  8'd10, 9'd284},{1'b0,  8'd11, 9'd198},{1'b0,  8'd14, 9'd323},{1'b0,  8'd18,  9'd56},{1'b0,  8'd28,   9'd0},{1'b0,  8'd35,  9'd77},{1'b0,  8'd48, 9'd188},{1'b0,  8'd58,   9'd0},{1'b0,  8'd74, 9'd295},{1'b0,  8'd85, 9'd233},{1'b0,  8'd88,   9'd0},{1'b0,  8'd92,  9'd10},{1'b0, 8'd110, 9'd298},{1'b0, 8'd118,   9'd0},{1'b0, 8'd127, 9'd254},{1'b1, 8'd128, 9'd182},
{1'b0,   8'd0, 9'd296},{1'b0,   8'd2,  9'd72},{1'b0,   8'd4,  9'd10},{1'b0,   8'd6, 9'd197},{1'b0,  8'd11, 9'd242},{1'b0,  8'd16, 9'd306},{1'b0,  8'd24,  9'd64},{1'b0,  8'd29,   9'd0},{1'b0,  8'd44,  9'd51},{1'b0,  8'd49, 9'd114},{1'b0,  8'd59,   9'd0},{1'b0,  8'd66, 9'd324},{1'b0,  8'd88, 9'd268},{1'b0,  8'd89,   9'd0},{1'b0,  8'd93,  9'd73},{1'b0,  8'd93, 9'd309},{1'b0, 8'd119,   9'd0},{1'b0, 8'd120,  9'd58},{1'b1, 8'd125, 9'd188}
};
localparam int          cLARGE_HS_TAB_8BY9_PACKED_SIZE = 500;
localparam bit [17 : 0] cLARGE_HS_TAB_8BY9_PACKED[cLARGE_HS_TAB_8BY9_PACKED_SIZE] = '{
{1'b0,   8'd0,   9'd0},{1'b0,   8'd1, 9'd290},{1'b0,  8'd15, 9'd196},{1'b0,  8'd17, 9'd231},{1'b0,  8'd20,   9'd0},{1'b0,  8'd25, 9'd312},{1'b0,  8'd34, 9'd121},{1'b0,  8'd40,   9'd0},{1'b0,  8'd50,  9'd37},{1'b0,  8'd57, 9'd238},{1'b0,  8'd60,   9'd0},{1'b0,  8'd77,  9'd30},{1'b0,  8'd79,  9'd63},{1'b0,  8'd80,   9'd0},{1'b0,  8'd83,  9'd22},{1'b0,  8'd91, 9'd336},{1'b0, 8'd100,   9'd0},{1'b0, 8'd109, 9'd206},{1'b0, 8'd109, 9'd214},{1'b0, 8'd120,   9'd0},{1'b0, 8'd121, 9'd348},{1'b0, 8'd136, 9'd216},{1'b0, 8'd140,   9'd0},{1'b0, 8'd152,  9'd80},{1'b1, 8'd153,  9'd34},
{1'b0,   8'd1,   9'd0},{1'b0,   8'd3, 9'd348},{1'b0,   8'd8, 9'd188},{1'b0,  8'd17, 9'd119},{1'b0,  8'd21,   9'd0},{1'b0,  8'd30, 9'd328},{1'b0,  8'd35,  9'd49},{1'b0,  8'd41,   9'd0},{1'b0,  8'd43,  9'd80},{1'b0,  8'd59, 9'd307},{1'b0,  8'd61,   9'd0},{1'b0,  8'd63,  9'd53},{1'b0,  8'd66, 9'd291},{1'b0,  8'd81,   9'd0},{1'b0,  8'd86,  9'd74},{1'b0,  8'd92, 9'd226},{1'b0, 8'd101,   9'd0},{1'b0, 8'd108, 9'd112},{1'b0, 8'd115, 9'd330},{1'b0, 8'd121,   9'd0},{1'b0, 8'd136, 9'd306},{1'b0, 8'd137, 9'd198},{1'b0, 8'd141,   9'd0},{1'b0, 8'd154,  9'd90},{1'b1, 8'd156,  9'd84},
{1'b0,   8'd0, 9'd161},{1'b0,   8'd2,   9'd0},{1'b0,   8'd7, 9'd317},{1'b0,  8'd17,  9'd74},{1'b0,  8'd22,   9'd0},{1'b0,  8'd29, 9'd261},{1'b0,  8'd38, 9'd190},{1'b0,  8'd42,   9'd0},{1'b0,  8'd43, 9'd281},{1'b0,  8'd55, 9'd235},{1'b0,  8'd62,   9'd0},{1'b0,  8'd72, 9'd349},{1'b0,  8'd76, 9'd242},{1'b0,  8'd82,   9'd0},{1'b0,  8'd91, 9'd181},{1'b0,  8'd98,  9'd88},{1'b0, 8'd101, 9'd103},{1'b0, 8'd102,   9'd0},{1'b0, 8'd105, 9'd118},{1'b0, 8'd122,   9'd0},{1'b0, 8'd122, 9'd353},{1'b0, 8'd128, 9'd123},{1'b0, 8'd142,   9'd0},{1'b0, 8'd148, 9'd260},{1'b1, 8'd149, 9'd236},
{1'b0,   8'd3,   9'd0},{1'b0,   8'd5, 9'd184},{1'b0,  8'd13,  9'd67},{1'b0,  8'd13, 9'd296},{1'b0,  8'd23,   9'd0},{1'b0,  8'd26, 9'd117},{1'b0,  8'd36, 9'd208},{1'b0,  8'd43,   9'd0},{1'b0,  8'd45, 9'd289},{1'b0,  8'd53, 9'd112},{1'b0,  8'd63,   9'd0},{1'b0,  8'd63, 9'd173},{1'b0,  8'd79, 9'd245},{1'b0,  8'd82,  9'd29},{1'b0,  8'd83,   9'd0},{1'b0,  8'd90, 9'd200},{1'b0, 8'd103,   9'd0},{1'b0, 8'd114,  9'd70},{1'b0, 8'd115, 9'd259},{1'b0, 8'd123,   9'd0},{1'b0, 8'd131, 9'd312},{1'b0, 8'd134, 9'd173},{1'b0, 8'd143,   9'd0},{1'b0, 8'd145, 9'd202},{1'b1, 8'd156, 9'd123},
{1'b0,   8'd4,   9'd0},{1'b0,   8'd4, 9'd313},{1'b0,   8'd9,  9'd13},{1'b0,  8'd16,  9'd82},{1'b0,  8'd21,  9'd75},{1'b0,  8'd22,  9'd95},{1'b0,  8'd24,   9'd0},{1'b0,  8'd44,   9'd0},{1'b0,  8'd44,  9'd26},{1'b0,  8'd51, 9'd147},{1'b0,  8'd64,   9'd0},{1'b0,  8'd71, 9'd179},{1'b0,  8'd74, 9'd248},{1'b0,  8'd81, 9'd161},{1'b0,  8'd84,   9'd0},{1'b0,  8'd93,  9'd58},{1'b0, 8'd104,   9'd0},{1'b0, 8'd118, 9'd309},{1'b0, 8'd119, 9'd338},{1'b0, 8'd123, 9'd180},{1'b0, 8'd124,   9'd0},{1'b0, 8'd132, 9'd132},{1'b0, 8'd144,   9'd0},{1'b0, 8'd149, 9'd151},{1'b1, 8'd158, 9'd214},
{1'b0,   8'd5,   9'd0},{1'b0,   8'd5, 9'd121},{1'b0,  8'd12, 9'd243},{1'b0,  8'd12, 9'd300},{1'b0,  8'd25,   9'd0},{1'b0,  8'd27, 9'd273},{1'b0,  8'd31, 9'd238},{1'b0,  8'd44, 9'd300},{1'b0,  8'd45,   9'd0},{1'b0,  8'd56, 9'd114},{1'b0,  8'd61,   9'd7},{1'b0,  8'd65,   9'd0},{1'b0,  8'd76, 9'd246},{1'b0,  8'd85,   9'd0},{1'b0,  8'd89, 9'd103},{1'b0,  8'd94,  9'd98},{1'b0, 8'd105,   9'd0},{1'b0, 8'd110, 9'd291},{1'b0, 8'd114,  9'd16},{1'b0, 8'd125,   9'd0},{1'b0, 8'd127, 9'd125},{1'b0, 8'd137,  9'd56},{1'b0, 8'd144, 9'd194},{1'b0, 8'd145,   9'd0},{1'b1, 8'd150, 9'd272},
{1'b0,   8'd6,   9'd0},{1'b0,   8'd9, 9'd145},{1'b0,  8'd12, 9'd164},{1'b0,  8'd19, 9'd189},{1'b0,  8'd20, 9'd308},{1'b0,  8'd26,   9'd0},{1'b0,  8'd32, 9'd298},{1'b0,  8'd40, 9'd306},{1'b0,  8'd46,   9'd0},{1'b0,  8'd49, 9'd128},{1'b0,  8'd60, 9'd253},{1'b0,  8'd61,  9'd65},{1'b0,  8'd66,   9'd0},{1'b0,  8'd84, 9'd311},{1'b0,  8'd86,   9'd0},{1'b0,  8'd95,   9'd3},{1'b0, 8'd106,   9'd0},{1'b0, 8'd106,  9'd61},{1'b0, 8'd117, 9'd242},{1'b0, 8'd126,   9'd0},{1'b0, 8'd128, 9'd240},{1'b0, 8'd135, 9'd265},{1'b0, 8'd143, 9'd311},{1'b0, 8'd144,  9'd72},{1'b1, 8'd146,   9'd0},
{1'b0,   8'd2,  9'd46},{1'b0,   8'd5,  9'd96},{1'b0,   8'd7,   9'd0},{1'b0,   8'd9, 9'd296},{1'b0,  8'd23, 9'd301},{1'b0,  8'd23, 9'd159},{1'b0,  8'd27,   9'd0},{1'b0,  8'd47,   9'd0},{1'b0,  8'd54,  9'd43},{1'b0,  8'd59, 9'd176},{1'b0,  8'd64, 9'd332},{1'b0,  8'd67,   9'd0},{1'b0,  8'd70,  9'd50},{1'b0,  8'd86, 9'd342},{1'b0,  8'd87,   9'd0},{1'b0,  8'd88, 9'd105},{1'b0, 8'd107,   9'd0},{1'b0, 8'd113, 9'd285},{1'b0, 8'd119, 9'd356},{1'b0, 8'd127,   9'd0},{1'b0, 8'd127, 9'd170},{1'b0, 8'd131, 9'd331},{1'b0, 8'd141, 9'd329},{1'b0, 8'd145, 9'd195},{1'b1, 8'd147,   9'd0},
{1'b0,   8'd0, 9'd142},{1'b0,   8'd1, 9'd267},{1'b0,   8'd8,   9'd0},{1'b0,   8'd8, 9'd121},{1'b0,  8'd28,   9'd0},{1'b0,  8'd29,  9'd79},{1'b0,  8'd39, 9'd197},{1'b0,  8'd48,   9'd0},{1'b0,  8'd51,  9'd97},{1'b0,  8'd52, 9'd326},{1'b0,  8'd60, 9'd107},{1'b0,  8'd68,   9'd0},{1'b0,  8'd70, 9'd246},{1'b0,  8'd82, 9'd151},{1'b0,  8'd88,   9'd0},{1'b0,  8'd90, 9'd319},{1'b0, 8'd103,  9'd61},{1'b0, 8'd107, 9'd227},{1'b0, 8'd108,   9'd0},{1'b0, 8'd128,   9'd0},{1'b0, 8'd130, 9'd267},{1'b0, 8'd133, 9'd254},{1'b0, 8'd148,   9'd0},{1'b0, 8'd151,  9'd91},{1'b1, 8'd158, 9'd286},
{1'b0,   8'd6, 9'd315},{1'b0,   8'd9,   9'd0},{1'b0,  8'd13, 9'd176},{1'b0,  8'd14, 9'd229},{1'b0,  8'd29,   9'd0},{1'b0,  8'd33,  9'd98},{1'b0,  8'd33, 9'd193},{1'b0,  8'd41,  9'd95},{1'b0,  8'd49,   9'd0},{1'b0,  8'd50,  9'd62},{1'b0,  8'd69,   9'd0},{1'b0,  8'd72, 9'd143},{1'b0,  8'd78, 9'd325},{1'b0,  8'd80, 9'd168},{1'b0,  8'd88,  9'd82},{1'b0,  8'd89,   9'd0},{1'b0, 8'd109,   9'd0},{1'b0, 8'd116, 9'd318},{1'b0, 8'd116, 9'd228},{1'b0, 8'd126, 9'd166},{1'b0, 8'd129,   9'd0},{1'b0, 8'd134, 9'd194},{1'b0, 8'd148, 9'd213},{1'b0, 8'd149,   9'd0},{1'b1, 8'd155, 9'd133},
{1'b0,   8'd2,   9'd4},{1'b0,   8'd7, 9'd153},{1'b0,  8'd10,   9'd0},{1'b0,  8'd10,  9'd97},{1'b0,  8'd22,   9'd6},{1'b0,  8'd25, 9'd143},{1'b0,  8'd30,   9'd0},{1'b0,  8'd42,  9'd42},{1'b0,  8'd49, 9'd171},{1'b0,  8'd50,   9'd0},{1'b0,  8'd68, 9'd196},{1'b0,  8'd70,   9'd0},{1'b0,  8'd75, 9'd220},{1'b0,  8'd90,   9'd0},{1'b0,  8'd93, 9'd352},{1'b0,  8'd96, 9'd148},{1'b0, 8'd100,  9'd48},{1'b0, 8'd102, 9'd243},{1'b0, 8'd110,   9'd0},{1'b0, 8'd122, 9'd135},{1'b0, 8'd125,   9'd5},{1'b0, 8'd130,   9'd0},{1'b0, 8'd150,   9'd0},{1'b0, 8'd151,  9'd18},{1'b1, 8'd154, 9'd334},
{1'b0,  8'd11,   9'd0},{1'b0,  8'd11, 9'd174},{1'b0,  8'd16,  9'd59},{1'b0,  8'd18, 9'd339},{1'b0,  8'd26,  9'd65},{1'b0,  8'd31,   9'd0},{1'b0,  8'd34, 9'd178},{1'b0,  8'd45, 9'd262},{1'b0,  8'd48,  9'd64},{1'b0,  8'd51,   9'd0},{1'b0,  8'd62,  9'd43},{1'b0,  8'd69,  9'd10},{1'b0,  8'd71,   9'd0},{1'b0,  8'd80, 9'd151},{1'b0,  8'd91,   9'd0},{1'b0,  8'd95, 9'd216},{1'b0, 8'd107, 9'd345},{1'b0, 8'd111,   9'd0},{1'b0, 8'd112, 9'd273},{1'b0, 8'd120,  9'd97},{1'b0, 8'd131,   9'd0},{1'b0, 8'd139, 9'd325},{1'b0, 8'd142,  9'd55},{1'b0, 8'd151,   9'd0},{1'b1, 8'd157, 9'd258},
{1'b0,   8'd1, 9'd174},{1'b0,   8'd4,  9'd58},{1'b0,  8'd12,   9'd0},{1'b0,  8'd14, 9'd106},{1'b0,  8'd32,   9'd0},{1'b0,  8'd32, 9'd344},{1'b0,  8'd35, 9'd231},{1'b0,  8'd46,   9'd8},{1'b0,  8'd46, 9'd101},{1'b0,  8'd52,   9'd0},{1'b0,  8'd66, 9'd246},{1'b0,  8'd72,   9'd0},{1'b0,  8'd73,  9'd80},{1'b0,  8'd87,  9'd96},{1'b0,  8'd92,   9'd0},{1'b0,  8'd97, 9'd232},{1'b0, 8'd100, 9'd128},{1'b0, 8'd112,   9'd0},{1'b0, 8'd118, 9'd354},{1'b0, 8'd132,   9'd0},{1'b0, 8'd133, 9'd210},{1'b0, 8'd139,  9'd39},{1'b0, 8'd150, 9'd318},{1'b0, 8'd152,   9'd0},{1'b1, 8'd157, 9'd298},
{1'b0,   8'd8,  9'd30},{1'b0,  8'd10, 9'd213},{1'b0,  8'd11, 9'd230},{1'b0,  8'd13,   9'd0},{1'b0,  8'd28, 9'd125},{1'b0,  8'd33,   9'd0},{1'b0,  8'd37,  9'd48},{1'b0,  8'd41,  9'd28},{1'b0,  8'd53,   9'd0},{1'b0,  8'd54, 9'd186},{1'b0,  8'd73,   9'd0},{1'b0,  8'd73,  9'd50},{1'b0,  8'd74,  9'd47},{1'b0,  8'd87, 9'd221},{1'b0,  8'd93,   9'd0},{1'b0,  8'd94, 9'd180},{1'b0, 8'd103, 9'd345},{1'b0, 8'd112, 9'd189},{1'b0, 8'd113,   9'd0},{1'b0, 8'd123,  9'd56},{1'b0, 8'd132, 9'd253},{1'b0, 8'd133,   9'd0},{1'b0, 8'd146, 9'd143},{1'b0, 8'd147,  9'd86},{1'b1, 8'd153,   9'd0},
{1'b0,   8'd6, 9'd185},{1'b0,   8'd7, 9'd357},{1'b0,  8'd14,   9'd0},{1'b0,  8'd18, 9'd300},{1'b0,  8'd31, 9'd102},{1'b0,  8'd34,   9'd0},{1'b0,  8'd39, 9'd189},{1'b0,  8'd42, 9'd201},{1'b0,  8'd54,   9'd0},{1'b0,  8'd55,  9'd68},{1'b0,  8'd64, 9'd277},{1'b0,  8'd69, 9'd154},{1'b0,  8'd74,   9'd0},{1'b0,  8'd85,  9'd54},{1'b0,  8'd92, 9'd184},{1'b0,  8'd94,   9'd0},{1'b0, 8'd110,  9'd23},{1'b0, 8'd111, 9'd107},{1'b0, 8'd114,   9'd0},{1'b0, 8'd124, 9'd184},{1'b0, 8'd129,  9'd10},{1'b0, 8'd134,   9'd0},{1'b0, 8'd140, 9'd196},{1'b0, 8'd153, 9'd103},{1'b1, 8'd154,   9'd0},
{1'b0,   8'd0, 9'd311},{1'b0,   8'd6, 9'd124},{1'b0,  8'd14, 9'd201},{1'b0,  8'd15,   9'd0},{1'b0,  8'd30,  9'd26},{1'b0,  8'd35,   9'd0},{1'b0,  8'd36, 9'd160},{1'b0,  8'd47,  9'd93},{1'b0,  8'd47, 9'd123},{1'b0,  8'd55,   9'd0},{1'b0,  8'd71,  9'd61},{1'b0,  8'd75,   9'd0},{1'b0,  8'd75, 9'd227},{1'b0,  8'd84, 9'd332},{1'b0,  8'd85, 9'd244},{1'b0,  8'd95,   9'd0},{1'b0, 8'd106,  9'd19},{1'b0, 8'd113,  9'd79},{1'b0, 8'd115,   9'd0},{1'b0, 8'd125,  9'd67},{1'b0, 8'd135,   9'd0},{1'b0, 8'd138,  9'd59},{1'b0, 8'd147, 9'd280},{1'b0, 8'd152, 9'd234},{1'b1, 8'd155,   9'd0},
{1'b0,   8'd3, 9'd225},{1'b0,  8'd10,  9'd85},{1'b0,  8'd16,   9'd0},{1'b0,  8'd18, 9'd329},{1'b0,  8'd20, 9'd257},{1'b0,  8'd21, 9'd217},{1'b0,  8'd36,   9'd0},{1'b0,  8'd40, 9'd159},{1'b0,  8'd53, 9'd180},{1'b0,  8'd56,   9'd0},{1'b0,  8'd67, 9'd317},{1'b0,  8'd67, 9'd237},{1'b0,  8'd76,   9'd0},{1'b0,  8'd96,   9'd0},{1'b0,  8'd96,  9'd89},{1'b0,  8'd99, 9'd286},{1'b0, 8'd105, 9'd145},{1'b0, 8'd116,   9'd0},{1'b0, 8'd117,  9'd44},{1'b0, 8'd126, 9'd336},{1'b0, 8'd129, 9'd210},{1'b0, 8'd136,   9'd0},{1'b0, 8'd142, 9'd329},{1'b0, 8'd156,   9'd0},{1'b1, 8'd159,  9'd84},
{1'b0,   8'd2, 9'd137},{1'b0,   8'd4, 9'd161},{1'b0,  8'd15, 9'd336},{1'b0,  8'd17,   9'd0},{1'b0,  8'd28, 9'd330},{1'b0,  8'd37,   9'd0},{1'b0,  8'd37, 9'd155},{1'b0,  8'd48,  9'd24},{1'b0,  8'd57,   9'd0},{1'b0,  8'd57, 9'd195},{1'b0,  8'd65, 9'd291},{1'b0,  8'd77,   9'd0},{1'b0,  8'd78, 9'd120},{1'b0,  8'd81, 9'd177},{1'b0,  8'd97,   9'd0},{1'b0,  8'd98, 9'd238},{1'b0, 8'd102, 9'd229},{1'b0, 8'd104,  9'd51},{1'b0, 8'd117,   9'd0},{1'b0, 8'd121, 9'd155},{1'b0, 8'd124,  9'd32},{1'b0, 8'd137,   9'd0},{1'b0, 8'd143,  9'd72},{1'b0, 8'd155,  9'd68},{1'b1, 8'd157,   9'd0},
{1'b0,  8'd16, 9'd299},{1'b0,  8'd18,   9'd0},{1'b0,  8'd19, 9'd136},{1'b0,  8'd19, 9'd295},{1'b0,  8'd24, 9'd335},{1'b0,  8'd38,   9'd0},{1'b0,  8'd38, 9'd309},{1'b0,  8'd56, 9'd234},{1'b0,  8'd58,   9'd0},{1'b0,  8'd58, 9'd202},{1'b0,  8'd68,  9'd20},{1'b0,  8'd77, 9'd288},{1'b0,  8'd78,   9'd0},{1'b0,  8'd83, 9'd162},{1'b0,  8'd97, 9'd160},{1'b0,  8'd98,   9'd0},{1'b0, 8'd108, 9'd230},{1'b0, 8'd111, 9'd277},{1'b0, 8'd118,   9'd0},{1'b0, 8'd120, 9'd317},{1'b0, 8'd135,  9'd23},{1'b0, 8'd138,   9'd0},{1'b0, 8'd140, 9'd138},{1'b0, 8'd141, 9'd161},{1'b1, 8'd158,   9'd0},
{1'b0,   8'd3, 9'd236},{1'b0,  8'd11, 9'd308},{1'b0,  8'd15,  9'd78},{1'b0,  8'd19,   9'd0},{1'b0,  8'd24,  9'd37},{1'b0,  8'd27,  9'd51},{1'b0,  8'd39,   9'd0},{1'b0,  8'd52, 9'd144},{1'b0,  8'd58,  9'd92},{1'b0,  8'd59,   9'd0},{1'b0,  8'd62, 9'd115},{1'b0,  8'd65,  9'd16},{1'b0,  8'd79,   9'd0},{1'b0,  8'd89, 9'd105},{1'b0,  8'd99,   9'd0},{1'b0,  8'd99,  9'd69},{1'b0, 8'd101, 9'd329},{1'b0, 8'd104, 9'd207},{1'b0, 8'd119,   9'd0},{1'b0, 8'd130, 9'd280},{1'b0, 8'd138, 9'd284},{1'b0, 8'd139,   9'd0},{1'b0, 8'd146, 9'd341},{1'b0, 8'd159,   9'd0},{1'b1, 8'd159,  9'd72}
};
localparam int          cLARGE_HS_TAB_9BY10_PACKED_SIZE = 504;
localparam bit [17 : 0] cLARGE_HS_TAB_9BY10_PACKED[cLARGE_HS_TAB_9BY10_PACKED_SIZE] = '{
{1'b0,   8'd0,   9'd0},{1'b0,   8'd1, 9'd290},{1'b0,  8'd11, 9'd300},{1'b0,  8'd13, 9'd196},{1'b0,  8'd18,   9'd0},{1'b0,  8'd26, 9'd312},{1'b0,  8'd35, 9'd121},{1'b0,  8'd36,   9'd0},{1'b0,  8'd37, 9'd208},{1'b0,  8'd53, 9'd126},{1'b0,  8'd54,   9'd0},{1'b0,  8'd57, 9'd114},{1'b0,  8'd64, 9'd291},{1'b0,  8'd72,   9'd0},{1'b0,  8'd84,  9'd74},{1'b0,  8'd86, 9'd103},{1'b0,  8'd90,   9'd0},{1'b0,  8'd91,   9'd8},{1'b0,  8'd97, 9'd237},{1'b0, 8'd108,   9'd0},{1'b0, 8'd112, 9'd348},{1'b0, 8'd124, 9'd216},{1'b0, 8'd126,   9'd0},{1'b0, 8'd126,  9'd94},{1'b0, 8'd131,  9'd58},{1'b0, 8'd144,   9'd0},{1'b0, 8'd153,  9'd65},{1'b1, 8'd154,  9'd64},
{1'b0,   8'd1,   9'd0},{1'b0,   8'd3, 9'd348},{1'b0,   8'd7, 9'd188},{1'b0,  8'd12, 9'd296},{1'b0,  8'd19,   9'd0},{1'b0,  8'd30, 9'd261},{1'b0,  8'd31, 9'd328},{1'b0,  8'd37,   9'd0},{1'b0,  8'd44, 9'd281},{1'b0,  8'd44,  9'd80},{1'b0,  8'd55,   9'd0},{1'b0,  8'd56, 9'd235},{1'b0,  8'd62, 9'd173},{1'b0,  8'd73,   9'd0},{1'b0,  8'd75,  9'd30},{1'b0,  8'd87, 9'd200},{1'b0,  8'd91,   9'd0},{1'b0,  8'd94, 9'd103},{1'b0, 8'd100, 9'd214},{1'b0, 8'd109,   9'd0},{1'b0, 8'd118, 9'd296},{1'b0, 8'd119,  9'd36},{1'b0, 8'd127,   9'd0},{1'b0, 8'd140,  9'd36},{1'b0, 8'd143, 9'd234},{1'b0, 8'd144, 9'd321},{1'b0, 8'd145,   9'd0},{1'b1, 8'd158, 9'd300},
{1'b0,   8'd0, 9'd161},{1'b0,   8'd2,   9'd0},{1'b0,   8'd8,  9'd13},{1'b0,  8'd16,  9'd74},{1'b0,  8'd20,   9'd0},{1'b0,  8'd27, 9'd117},{1'b0,  8'd34, 9'd193},{1'b0,  8'd36,  9'd49},{1'b0,  8'd38,   9'd0},{1'b0,  8'd40, 9'd189},{1'b0,  8'd56,   9'd0},{1'b0,  8'd58, 9'd238},{1'b0,  8'd62,  9'd53},{1'b0,  8'd74,   9'd0},{1'b0,  8'd79, 9'd229},{1'b0,  8'd82, 9'd243},{1'b0,  8'd92,   9'd0},{1'b0,  8'd98, 9'd112},{1'b0, 8'd100, 9'd206},{1'b0, 8'd109, 9'd289},{1'b0, 8'd110,   9'd0},{1'b0, 8'd124, 9'd306},{1'b0, 8'd128,   9'd0},{1'b0, 8'd137, 9'd260},{1'b0, 8'd143,  9'd80},{1'b0, 8'd146,   9'd0},{1'b0, 8'd146,  9'd84},{1'b1, 8'd159, 9'd282},
{1'b0,   8'd3,   9'd0},{1'b0,   8'd5, 9'd184},{1'b0,  8'd12,  9'd67},{1'b0,  8'd16, 9'd119},{1'b0,  8'd20, 9'd189},{1'b0,  8'd21,   9'd0},{1'b0,  8'd23,  9'd95},{1'b0,  8'd39,   9'd0},{1'b0,  8'd39, 9'd190},{1'b0,  8'd52,  9'd37},{1'b0,  8'd57,   9'd0},{1'b0,  8'd69, 9'd179},{1'b0,  8'd71,  9'd50},{1'b0,  8'd75,   9'd0},{1'b0,  8'd78,  9'd29},{1'b0,  8'd79,  9'd60},{1'b0,  8'd93,   9'd0},{1'b0, 8'd105,  9'd70},{1'b0, 8'd106, 9'd259},{1'b0, 8'd108, 9'd176},{1'b0, 8'd110, 9'd309},{1'b0, 8'd111,   9'd0},{1'b0, 8'd129,   9'd0},{1'b0, 8'd135, 9'd202},{1'b0, 8'd138, 9'd169},{1'b0, 8'd146, 9'd123},{1'b0, 8'd147,   9'd0},{1'b1, 8'd152,  9'd75},
{1'b0,   8'd4,   9'd0},{1'b0,   8'd4, 9'd313},{1'b0,   8'd5, 9'd121},{1'b0,  8'd14,  9'd82},{1'b0,  8'd22,   9'd0},{1'b0,  8'd22,  9'd75},{1'b0,  8'd24, 9'd159},{1'b0,  8'd40,   9'd0},{1'b0,  8'd45,  9'd33},{1'b0,  8'd51, 9'd128},{1'b0,  8'd58,   9'd0},{1'b0,  8'd61,  9'd65},{1'b0,  8'd68, 9'd246},{1'b0,  8'd76,   9'd0},{1'b0,  8'd77, 9'd161},{1'b0,  8'd80, 9'd129},{1'b0,  8'd90,  9'd98},{1'b0,  8'd90, 9'd180},{1'b0,  8'd94,   9'd0},{1'b0, 8'd112,   9'd0},{1'b0, 8'd114, 9'd180},{1'b0, 8'd115, 9'd223},{1'b0, 8'd126, 9'd324},{1'b0, 8'd130,   9'd0},{1'b0, 8'd134, 9'd194},{1'b0, 8'd148,   9'd0},{1'b0, 8'd152, 9'd277},{1'b1, 8'd155, 9'd298},
{1'b0,   8'd5,   9'd0},{1'b0,   8'd8, 9'd145},{1'b0,  8'd11, 9'd164},{1'b0,  8'd16, 9'd231},{1'b0,  8'd18, 9'd300},{1'b0,  8'd23,   9'd0},{1'b0,  8'd32, 9'd238},{1'b0,  8'd41,   9'd0},{1'b0,  8'd46, 9'd300},{1'b0,  8'd46,  9'd26},{1'b0,  8'd59,   9'd0},{1'b0,  8'd59, 9'd307},{1'b0,  8'd61,   9'd7},{1'b0,  8'd74, 9'd246},{1'b0,  8'd74, 9'd242},{1'b0,  8'd77,   9'd0},{1'b0,  8'd92,  9'd88},{1'b0,  8'd95,   9'd0},{1'b0, 8'd105,  9'd16},{1'b0, 8'd113,   9'd0},{1'b0, 8'd121, 9'd211},{1'b0, 8'd122, 9'd173},{1'b0, 8'd131,   9'd0},{1'b0, 8'd132, 9'd351},{1'b0, 8'd133, 9'd311},{1'b0, 8'd149,   9'd0},{1'b0, 8'd149,  9'd84},{1'b1, 8'd159, 9'd149},
{1'b0,   8'd2,  9'd46},{1'b0,   8'd5,  9'd96},{1'b0,   8'd6,   9'd0},{1'b0,   8'd8, 9'd296},{1'b0,  8'd19, 9'd166},{1'b0,  8'd21, 9'd308},{1'b0,  8'd24,   9'd0},{1'b0,  8'd40, 9'd197},{1'b0,  8'd42,   9'd0},{1'b0,  8'd52,  9'd62},{1'b0,  8'd60,   9'd0},{1'b0,  8'd60, 9'd253},{1'b0,  8'd68,  9'd50},{1'b0,  8'd78,   9'd0},{1'b0,  8'd78, 9'd151},{1'b0,  8'd87, 9'd319},{1'b0,  8'd93, 9'd286},{1'b0,  8'd95, 9'd150},{1'b0,  8'd96,   9'd0},{1'b0, 8'd113, 9'd145},{1'b0, 8'd114,   9'd0},{1'b0, 8'd121, 9'd279},{1'b0, 8'd132,   9'd0},{1'b0, 8'd135, 9'd195},{1'b0, 8'd139, 9'd145},{1'b0, 8'd148, 9'd214},{1'b0, 8'd150,   9'd0},{1'b1, 8'd151, 9'd293},
{1'b0,   8'd0, 9'd142},{1'b0,   8'd1, 9'd267},{1'b0,   8'd7,   9'd0},{1'b0,   8'd7, 9'd121},{1'b0,  8'd24, 9'd301},{1'b0,  8'd25,   9'd0},{1'b0,  8'd28, 9'd273},{1'b0,  8'd36, 9'd231},{1'b0,  8'd41, 9'd306},{1'b0,  8'd43,   9'd0},{1'b0,  8'd56,  9'd68},{1'b0,  8'd58, 9'd195},{1'b0,  8'd61,   9'd0},{1'b0,  8'd79,   9'd0},{1'b0,  8'd81, 9'd311},{1'b0,  8'd84, 9'd342},{1'b0,  8'd91, 9'd119},{1'b0,  8'd92, 9'd238},{1'b0,  8'd97,   9'd0},{1'b0, 8'd115,   9'd0},{1'b0, 8'd116, 9'd125},{1'b0, 8'd116, 9'd170},{1'b0, 8'd133,   9'd0},{1'b0, 8'd134,  9'd72},{1'b0, 8'd136, 9'd127},{1'b0, 8'd148, 9'd286},{1'b0, 8'd151,   9'd0},{1'b1, 8'd156,  9'd78},
{1'b0,   8'd6, 9'd315},{1'b0,   8'd8,   9'd0},{1'b0,  8'd11, 9'd243},{1'b0,  8'd17,  9'd14},{1'b0,  8'd26,   9'd0},{1'b0,  8'd26, 9'd143},{1'b0,  8'd30,  9'd79},{1'b0,  8'd44,   9'd0},{1'b0,  8'd47, 9'd262},{1'b0,  8'd47, 9'd289},{1'b0,  8'd55,  9'd43},{1'b0,  8'd62,   9'd0},{1'b0,  8'd63,  9'd60},{1'b0,  8'd80,   9'd0},{1'b0,  8'd88, 9'd336},{1'b0,  8'd88, 9'd181},{1'b0,  8'd98,   9'd0},{1'b0, 8'd102, 9'd341},{1'b0, 8'd107, 9'd354},{1'b0, 8'd109, 9'd117},{1'b0, 8'd116,   9'd0},{1'b0, 8'd118,  9'd66},{1'b0, 8'd131,  9'd82},{1'b0, 8'd134,   9'd0},{1'b0, 8'd141, 9'd346},{1'b0, 8'd150, 9'd175},{1'b0, 8'd152,   9'd0},{1'b1, 8'd161, 9'd188},
{1'b0,   8'd2,   9'd4},{1'b0,   8'd9,   9'd0},{1'b0,   8'd9,  9'd97},{1'b0,  8'd15, 9'd213},{1'b0,  8'd23,   9'd6},{1'b0,  8'd27,   9'd0},{1'b0,  8'd27,  9'd65},{1'b0,  8'd42,  9'd95},{1'b0,  8'd43,  9'd42},{1'b0,  8'd45,   9'd0},{1'b0,  8'd60, 9'd107},{1'b0,  8'd63,   9'd0},{1'b0,  8'd70, 9'd143},{1'b0,  8'd72,  9'd47},{1'b0,  8'd80, 9'd333},{1'b0,  8'd81,   9'd0},{1'b0,  8'd97,  9'd38},{1'b0,  8'd99,   9'd0},{1'b0, 8'd106, 9'd330},{1'b0, 8'd117,   9'd0},{1'b0, 8'd120, 9'd254},{1'b0, 8'd123, 9'd265},{1'b0, 8'd128, 9'd342},{1'b0, 8'd135,   9'd0},{1'b0, 8'd140, 9'd181},{1'b0, 8'd145, 9'd133},{1'b0, 8'd153,   9'd0},{1'b1, 8'd160,  9'd97},
{1'b0,  8'd10,   9'd0},{1'b0,  8'd10, 9'd174},{1'b0,  8'd14,  9'd59},{1'b0,  8'd17, 9'd131},{1'b0,  8'd28,   9'd0},{1'b0,  8'd32, 9'd102},{1'b0,  8'd33, 9'd298},{1'b0,  8'd38,  9'd48},{1'b0,  8'd46,   9'd0},{1'b0,  8'd51, 9'd171},{1'b0,  8'd54, 9'd326},{1'b0,  8'd64,   9'd0},{1'b0,  8'd67, 9'd154},{1'b0,  8'd73, 9'd220},{1'b0,  8'd82,   9'd0},{1'b0,  8'd89, 9'd184},{1'b0,  8'd93,  9'd69},{1'b0, 8'd100,   9'd0},{1'b0, 8'd104, 9'd285},{1'b0, 8'd108, 9'd260},{1'b0, 8'd114,  9'd56},{1'b0, 8'd118,   9'd0},{1'b0, 8'd132, 9'd224},{1'b0, 8'd136,   9'd0},{1'b0, 8'd139, 9'd156},{1'b0, 8'd154,   9'd0},{1'b0, 8'd154, 9'd242},{1'b1, 8'd160,  9'd17},
{1'b0,   8'd1, 9'd174},{1'b0,   8'd4,  9'd58},{1'b0,  8'd11,   9'd0},{1'b0,  8'd12, 9'd176},{1'b0,  8'd29,   9'd0},{1'b0,  8'd29, 9'd125},{1'b0,  8'd34,  9'd98},{1'b0,  8'd38, 9'd155},{1'b0,  8'd47,   9'd0},{1'b0,  8'd48,   9'd8},{1'b0,  8'd55, 9'd186},{1'b0,  8'd65,   9'd0},{1'b0,  8'd67,  9'd10},{1'b0,  8'd72, 9'd248},{1'b0,  8'd73, 9'd227},{1'b0,  8'd83,   9'd0},{1'b0, 8'd101,   9'd0},{1'b0, 8'd101, 9'd284},{1'b0, 8'd102, 9'd184},{1'b0, 8'd111,  9'd97},{1'b0, 8'd119,   9'd0},{1'b0, 8'd120, 9'd210},{1'b0, 8'd130, 9'd123},{1'b0, 8'd137,   9'd0},{1'b0, 8'd137, 9'd213},{1'b0, 8'd147, 9'd311},{1'b0, 8'd155,   9'd0},{1'b1, 8'd161, 9'd110},
{1'b0,   8'd6, 9'd185},{1'b0,   8'd7,  9'd30},{1'b0,   8'd9, 9'd213},{1'b0,  8'd12,   9'd0},{1'b0,  8'd30,   9'd0},{1'b0,  8'd31,  9'd26},{1'b0,  8'd35, 9'd178},{1'b0,  8'd42,  9'd28},{1'b0,  8'd48,   9'd0},{1'b0,  8'd50,  9'd64},{1'b0,  8'd64, 9'd246},{1'b0,  8'd66,   9'd0},{1'b0,  8'd66, 9'd196},{1'b0,  8'd76,  9'd63},{1'b0,  8'd83,  9'd54},{1'b0,  8'd84,   9'd0},{1'b0,  8'd96, 9'd186},{1'b0, 8'd102,   9'd0},{1'b0, 8'd107, 9'd252},{1'b0, 8'd110, 9'd354},{1'b0, 8'd119, 9'd217},{1'b0, 8'd120,   9'd0},{1'b0, 8'd129, 9'd196},{1'b0, 8'd130, 9'd352},{1'b0, 8'd138,   9'd0},{1'b0, 8'd144,  9'd88},{1'b0, 8'd156,   9'd0},{1'b1, 8'd158,  9'd85},
{1'b0,   8'd0, 9'd311},{1'b0,  8'd13,   9'd0},{1'b0,  8'd15,  9'd98},{1'b0,  8'd15, 9'd242},{1'b0,  8'd20,  9'd92},{1'b0,  8'd29, 9'd330},{1'b0,  8'd31,   9'd0},{1'b0,  8'd43, 9'd201},{1'b0,  8'd45, 9'd312},{1'b0,  8'd49,   9'd0},{1'b0,  8'd57, 9'd234},{1'b0,  8'd67,   9'd0},{1'b0,  8'd69,  9'd61},{1'b0,  8'd82,  9'd87},{1'b0,  8'd85,   9'd0},{1'b0,  8'd85, 9'd297},{1'b0, 8'd101,  9'd51},{1'b0, 8'd103,   9'd0},{1'b0, 8'd103, 9'd107},{1'b0, 8'd117, 9'd170},{1'b0, 8'd121,   9'd0},{1'b0, 8'd125, 9'd243},{1'b0, 8'd136, 9'd286},{1'b0, 8'd138,  9'd35},{1'b0, 8'd139,   9'd0},{1'b0, 8'd145,  9'd68},{1'b0, 8'd157,   9'd0},{1'b1, 8'd157, 9'd313},
{1'b0,   8'd3, 9'd225},{1'b0,   8'd6, 9'd124},{1'b0,  8'd10, 9'd230},{1'b0,  8'd14,   9'd0},{1'b0,  8'd19, 9'd242},{1'b0,  8'd21, 9'd257},{1'b0,  8'd32,   9'd0},{1'b0,  8'd41, 9'd159},{1'b0,  8'd48, 9'd101},{1'b0,  8'd50,   9'd0},{1'b0,  8'd65, 9'd237},{1'b0,  8'd68,   9'd0},{1'b0,  8'd70, 9'd349},{1'b0,  8'd75, 9'd288},{1'b0,  8'd81, 9'd332},{1'b0,  8'd86,   9'd0},{1'b0,  8'd95, 9'd267},{1'b0,  8'd99,  9'd41},{1'b0, 8'd104,   9'd0},{1'b0, 8'd113,  9'd66},{1'b0, 8'd122,   9'd0},{1'b0, 8'd122, 9'd194},{1'b0, 8'd127, 9'd284},{1'b0, 8'd140,   9'd0},{1'b0, 8'd142, 9'd163},{1'b0, 8'd147,  9'd39},{1'b0, 8'd153, 9'd313},{1'b1, 8'd158,   9'd0},
{1'b0,   8'd2, 9'd137},{1'b0,  8'd13, 9'd336},{1'b0,  8'd15,   9'd0},{1'b0,  8'd17, 9'd280},{1'b0,  8'd22, 9'd217},{1'b0,  8'd28,  9'd51},{1'b0,  8'd33,   9'd0},{1'b0,  8'd49,  9'd93},{1'b0,  8'd49, 9'd123},{1'b0,  8'd51,   9'd0},{1'b0,  8'd63, 9'd173},{1'b0,  8'd66,  9'd20},{1'b0,  8'd69,   9'd0},{1'b0,  8'd83, 9'd244},{1'b0,  8'd85, 9'd220},{1'b0,  8'd87,   9'd0},{1'b0,  8'd99, 9'd116},{1'b0, 8'd104,  9'd79},{1'b0, 8'd105,   9'd0},{1'b0, 8'd112, 9'd155},{1'b0, 8'd115, 9'd293},{1'b0, 8'd123,   9'd0},{1'b0, 8'd128, 9'd317},{1'b0, 8'd129, 9'd138},{1'b0, 8'd141,   9'd0},{1'b0, 8'd151, 9'd146},{1'b0, 8'd155, 9'd197},{1'b1, 8'd159,   9'd0},
{1'b0,   8'd4, 9'd161},{1'b0,   8'd9,  9'd85},{1'b0,  8'd14, 9'd299},{1'b0,  8'd16,   9'd0},{1'b0,  8'd18, 9'd339},{1'b0,  8'd33, 9'd344},{1'b0,  8'd34,   9'd0},{1'b0,  8'd37, 9'd160},{1'b0,  8'd52,   9'd0},{1'b0,  8'd53, 9'd319},{1'b0,  8'd59, 9'd176},{1'b0,  8'd65, 9'd317},{1'b0,  8'd70,   9'd0},{1'b0,  8'd76, 9'd245},{1'b0,  8'd77, 9'd177},{1'b0,  8'd88,   9'd0},{1'b0,  8'd98, 9'd230},{1'b0, 8'd103, 9'd277},{1'b0, 8'd106,   9'd0},{1'b0, 8'd111, 9'd317},{1'b0, 8'd124,   9'd0},{1'b0, 8'd125, 9'd226},{1'b0, 8'd127,  9'd59},{1'b0, 8'd142,   9'd0},{1'b0, 8'd142,  9'd35},{1'b0, 8'd149,  9'd72},{1'b0, 8'd150, 9'd141},{1'b1, 8'd160,   9'd0},
{1'b0,   8'd3, 9'd236},{1'b0,  8'd10, 9'd308},{1'b0,  8'd13,  9'd78},{1'b0,  8'd17,   9'd0},{1'b0,  8'd25, 9'd335},{1'b0,  8'd25,  9'd37},{1'b0,  8'd35,   9'd0},{1'b0,  8'd39, 9'd309},{1'b0,  8'd50,  9'd24},{1'b0,  8'd53,   9'd0},{1'b0,  8'd54, 9'd144},{1'b0,  8'd71,   9'd0},{1'b0,  8'd71,  9'd80},{1'b0,  8'd86, 9'd105},{1'b0,  8'd89,   9'd0},{1'b0,  8'd89, 9'd226},{1'b0,  8'd94, 9'd329},{1'b0,  8'd96,  9'd81},{1'b0, 8'd107,   9'd0},{1'b0, 8'd117, 9'd137},{1'b0, 8'd123,  9'd23},{1'b0, 8'd125,   9'd0},{1'b0, 8'd133,  9'd72},{1'b0, 8'd141,  9'd32},{1'b0, 8'd143,   9'd0},{1'b0, 8'd156, 9'd198},{1'b0, 8'd157, 9'd258},{1'b1, 8'd161,   9'd0}
};
