//
// Project       : rsc2
// Author        : Shekhalev Denis (des00)
// Workfile      : rsc2_dvb_ptable.svh
// Description   : file with RSC2 reordered permutation tables A-1/2/4/5
//

  localparam int cDVB_PTABLE_SIZE = 34;

  typedef int   tab_t     [6];  // {P, Q0, Q1, Q2, Q3, N}
  typedef tab_t tab_dvb_t [cDVB_PTABLE_SIZE];

  // {P, Q0, Q1, Q2, Q3, N}
  localparam tab_dvb_t cDVB_PTABLE = '{
    '{  9,   2,   2,   8,  0,  14 * 4 } , // 0
    '{ 17,   9,   5,  14,  1,  38 * 4 } , // 1
    '{ 23,  10,   5,   0,  0,  51 * 4 } , // 2
    '{ 23,   6,  10,   4,  0,  55 * 4 } , // 3
    '{ 23,  10,   2,  11,  1,  59 * 4 } , // 4
    '{ 23,   6,   8,   1,  1,  62 * 4 } , // 5
    '{ 25,   1,   1,   2,  0,  69 * 4 } , // 6
    '{ 23,   8,   1,   4,  1,  84 * 4 } , // 7
    '{ 23,   6,  13,  10,  0,  85 * 4 } , // 8
    '{ 25,   1,   7,   2,  1,  93 * 4 } , // 9
    '{ 25,   1,   2,   0,  1,  96 * 4 } , // 10
    '{ 23,  10,   8,   2,  1, 100 * 4 } , // 11
    '{ 29,   1,   4,   1,  1, 108 * 4 } , // 12
    '{ 29,   6,   5,   0,  0, 115 * 4 } , // 13
    '{ 31,   0,   3,   1,  0, 123 * 4 } , // 14
    '{ 31,   1,   1,   2,  1, 128 * 4 } , // 15
    '{ 31,   0,   1,   2,  0, 130 * 4 } , // 16
    '{ 31,   0,   0,   0,  0, 144 * 4 } , // 17
    '{ 33,   9,  15,   3,  1, 170 * 4 } , // 18
    '{ 37,   0,   2,   0,  2, 175 * 4 } , // 19
    '{ 37,   1,   3,   4,  2, 188 * 4 } , // 20
    '{ 37,   6,   1,  15,  0, 192 * 4 } , // 21
    '{ 39,   7,   0,   0,  0, 194 * 4 } , // 22
    '{ 45,   1,   1,   4,  0, 256 * 4 } , // 23
    '{ 43,   0,   0,   6,  2, 264 * 4 } , // 24
    '{ 49,   0,   3,   5,  0, 298 * 4 } , // 25
    '{ 49,   0,   6,   0,  1, 307 * 4 } , // 26
    '{ 49,   0,   5,   0,  5, 333 * 4 } , // 27
    '{ 53,   1,   4,   6,  2, 355 * 4 } , // 28
    '{ 53,   1,  10,   7,  1, 400 * 4 } , // 29
    '{ 59,   1,   1,   2,  1, 438 * 4 } , // 30
    '{ 59,   3,   8,   5,  1, 444 * 4 } , // 31
    '{ 65,   0,   3,   7,  0, 539 * 4 } , // 32
    '{ 81,   1,   2,   5,  2, 599 * 4 }   // 33
  };
